
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"cc",x"cf",x"c4",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"cc",x"cf",x"c4"),
    14 => (x"48",x"ec",x"ef",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e6",x"e7"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"4a",x"71",x"86",x"fc"),
    21 => (x"69",x"49",x"c0",x"ff"),
    22 => (x"98",x"c0",x"c4",x"48"),
    23 => (x"02",x"6e",x"7e",x"70"),
    24 => (x"79",x"72",x"87",x"f5"),
    25 => (x"26",x"8e",x"fc",x"48"),
    26 => (x"5b",x"5e",x"0e",x"4f"),
    27 => (x"4b",x"71",x"0e",x"5c"),
    28 => (x"4a",x"13",x"4c",x"c0"),
    29 => (x"87",x"cd",x"02",x"9a"),
    30 => (x"d2",x"ff",x"49",x"72"),
    31 => (x"13",x"84",x"c1",x"87"),
    32 => (x"f3",x"05",x"9a",x"4a"),
    33 => (x"26",x"48",x"74",x"87"),
    34 => (x"26",x"4b",x"26",x"4c"),
    35 => (x"1e",x"72",x"1e",x"4f"),
    36 => (x"48",x"12",x"1e",x"73"),
    37 => (x"87",x"ca",x"02",x"11"),
    38 => (x"98",x"df",x"c3",x"4b"),
    39 => (x"02",x"88",x"73",x"9b"),
    40 => (x"4b",x"26",x"87",x"f0"),
    41 => (x"4f",x"26",x"4a",x"26"),
    42 => (x"72",x"1e",x"73",x"1e"),
    43 => (x"04",x"8b",x"c1",x"1e"),
    44 => (x"48",x"12",x"87",x"ca"),
    45 => (x"87",x"c4",x"02",x"11"),
    46 => (x"87",x"f1",x"02",x"88"),
    47 => (x"4b",x"26",x"4a",x"26"),
    48 => (x"74",x"1e",x"4f",x"26"),
    49 => (x"72",x"1e",x"73",x"1e"),
    50 => (x"04",x"8b",x"c1",x"1e"),
    51 => (x"48",x"12",x"87",x"d0"),
    52 => (x"87",x"ca",x"02",x"11"),
    53 => (x"98",x"df",x"c3",x"4c"),
    54 => (x"02",x"88",x"74",x"9c"),
    55 => (x"4a",x"26",x"87",x"eb"),
    56 => (x"4c",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"a9",x"73",x"81",x"48"),
    59 => (x"12",x"87",x"c5",x"02"),
    60 => (x"87",x"f6",x"05",x"53"),
    61 => (x"c4",x"1e",x"4f",x"26"),
    62 => (x"48",x"71",x"4a",x"66"),
    63 => (x"fb",x"05",x"51",x"12"),
    64 => (x"1e",x"4f",x"26",x"87"),
    65 => (x"73",x"81",x"48",x"73"),
    66 => (x"53",x"72",x"05",x"a9"),
    67 => (x"4f",x"26",x"87",x"f9"),
    68 => (x"72",x"1e",x"73",x"1e"),
    69 => (x"e7",x"c0",x"02",x"9a"),
    70 => (x"c1",x"48",x"c0",x"87"),
    71 => (x"06",x"a9",x"72",x"4b"),
    72 => (x"82",x"72",x"87",x"d1"),
    73 => (x"73",x"87",x"c9",x"06"),
    74 => (x"01",x"a9",x"72",x"83"),
    75 => (x"87",x"c3",x"87",x"f4"),
    76 => (x"72",x"3a",x"b2",x"c1"),
    77 => (x"73",x"89",x"03",x"a9"),
    78 => (x"2a",x"c1",x"07",x"80"),
    79 => (x"87",x"f3",x"05",x"2b"),
    80 => (x"4f",x"26",x"4b",x"26"),
    81 => (x"c4",x"1e",x"75",x"1e"),
    82 => (x"a1",x"b7",x"71",x"4d"),
    83 => (x"c1",x"b9",x"ff",x"04"),
    84 => (x"07",x"bd",x"c3",x"81"),
    85 => (x"04",x"a2",x"b7",x"72"),
    86 => (x"82",x"c1",x"ba",x"ff"),
    87 => (x"fe",x"07",x"bd",x"c1"),
    88 => (x"2d",x"c1",x"87",x"ee"),
    89 => (x"c1",x"b8",x"ff",x"04"),
    90 => (x"04",x"2d",x"07",x"80"),
    91 => (x"81",x"c1",x"b9",x"ff"),
    92 => (x"26",x"4d",x"26",x"07"),
    93 => (x"48",x"11",x"1e",x"4f"),
    94 => (x"78",x"08",x"d4",x"ff"),
    95 => (x"c1",x"48",x"66",x"c4"),
    96 => (x"58",x"a6",x"c8",x"88"),
    97 => (x"ed",x"05",x"98",x"70"),
    98 => (x"1e",x"4f",x"26",x"87"),
    99 => (x"c3",x"48",x"d4",x"ff"),
   100 => (x"51",x"68",x"78",x"ff"),
   101 => (x"c1",x"48",x"66",x"c4"),
   102 => (x"58",x"a6",x"c8",x"88"),
   103 => (x"eb",x"05",x"98",x"70"),
   104 => (x"1e",x"4f",x"26",x"87"),
   105 => (x"d4",x"ff",x"1e",x"73"),
   106 => (x"7b",x"ff",x"c3",x"4b"),
   107 => (x"ff",x"c3",x"4a",x"6b"),
   108 => (x"c8",x"49",x"6b",x"7b"),
   109 => (x"c3",x"b1",x"72",x"32"),
   110 => (x"4a",x"6b",x"7b",x"ff"),
   111 => (x"b2",x"71",x"31",x"c8"),
   112 => (x"6b",x"7b",x"ff",x"c3"),
   113 => (x"72",x"32",x"c8",x"49"),
   114 => (x"c4",x"48",x"71",x"b1"),
   115 => (x"26",x"4d",x"26",x"87"),
   116 => (x"26",x"4b",x"26",x"4c"),
   117 => (x"5b",x"5e",x"0e",x"4f"),
   118 => (x"71",x"0e",x"5d",x"5c"),
   119 => (x"4c",x"d4",x"ff",x"4a"),
   120 => (x"ff",x"c3",x"49",x"72"),
   121 => (x"c3",x"7c",x"71",x"99"),
   122 => (x"05",x"bf",x"ec",x"ef"),
   123 => (x"66",x"d0",x"87",x"c8"),
   124 => (x"d4",x"30",x"c9",x"48"),
   125 => (x"66",x"d0",x"58",x"a6"),
   126 => (x"c3",x"29",x"d8",x"49"),
   127 => (x"7c",x"71",x"99",x"ff"),
   128 => (x"d0",x"49",x"66",x"d0"),
   129 => (x"99",x"ff",x"c3",x"29"),
   130 => (x"66",x"d0",x"7c",x"71"),
   131 => (x"c3",x"29",x"c8",x"49"),
   132 => (x"7c",x"71",x"99",x"ff"),
   133 => (x"c3",x"49",x"66",x"d0"),
   134 => (x"7c",x"71",x"99",x"ff"),
   135 => (x"29",x"d0",x"49",x"72"),
   136 => (x"71",x"99",x"ff",x"c3"),
   137 => (x"c9",x"4b",x"6c",x"7c"),
   138 => (x"c3",x"4d",x"ff",x"f0"),
   139 => (x"d0",x"05",x"ab",x"ff"),
   140 => (x"7c",x"ff",x"c3",x"87"),
   141 => (x"8d",x"c1",x"4b",x"6c"),
   142 => (x"c3",x"87",x"c6",x"02"),
   143 => (x"f0",x"02",x"ab",x"ff"),
   144 => (x"fe",x"48",x"73",x"87"),
   145 => (x"c0",x"1e",x"87",x"c7"),
   146 => (x"48",x"d4",x"ff",x"49"),
   147 => (x"c1",x"78",x"ff",x"c3"),
   148 => (x"b7",x"c8",x"c3",x"81"),
   149 => (x"87",x"f1",x"04",x"a9"),
   150 => (x"73",x"1e",x"4f",x"26"),
   151 => (x"c4",x"87",x"e7",x"1e"),
   152 => (x"c0",x"4b",x"df",x"f8"),
   153 => (x"f0",x"ff",x"c0",x"1e"),
   154 => (x"fd",x"49",x"f7",x"c1"),
   155 => (x"86",x"c4",x"87",x"e7"),
   156 => (x"c0",x"05",x"a8",x"c1"),
   157 => (x"d4",x"ff",x"87",x"ea"),
   158 => (x"78",x"ff",x"c3",x"48"),
   159 => (x"c0",x"c0",x"c0",x"c1"),
   160 => (x"c0",x"1e",x"c0",x"c0"),
   161 => (x"e9",x"c1",x"f0",x"e1"),
   162 => (x"87",x"c9",x"fd",x"49"),
   163 => (x"98",x"70",x"86",x"c4"),
   164 => (x"ff",x"87",x"ca",x"05"),
   165 => (x"ff",x"c3",x"48",x"d4"),
   166 => (x"cb",x"48",x"c1",x"78"),
   167 => (x"87",x"e6",x"fe",x"87"),
   168 => (x"fe",x"05",x"8b",x"c1"),
   169 => (x"48",x"c0",x"87",x"fd"),
   170 => (x"1e",x"87",x"e6",x"fc"),
   171 => (x"d4",x"ff",x"1e",x"73"),
   172 => (x"78",x"ff",x"c3",x"48"),
   173 => (x"1e",x"c0",x"4b",x"d3"),
   174 => (x"c1",x"f0",x"ff",x"c0"),
   175 => (x"d4",x"fc",x"49",x"c1"),
   176 => (x"70",x"86",x"c4",x"87"),
   177 => (x"87",x"ca",x"05",x"98"),
   178 => (x"c3",x"48",x"d4",x"ff"),
   179 => (x"48",x"c1",x"78",x"ff"),
   180 => (x"f1",x"fd",x"87",x"cb"),
   181 => (x"05",x"8b",x"c1",x"87"),
   182 => (x"c0",x"87",x"db",x"ff"),
   183 => (x"87",x"f1",x"fb",x"48"),
   184 => (x"5c",x"5b",x"5e",x"0e"),
   185 => (x"4c",x"d4",x"ff",x"0e"),
   186 => (x"c6",x"87",x"db",x"fd"),
   187 => (x"e1",x"c0",x"1e",x"ea"),
   188 => (x"49",x"c8",x"c1",x"f0"),
   189 => (x"c4",x"87",x"de",x"fb"),
   190 => (x"02",x"a8",x"c1",x"86"),
   191 => (x"ea",x"fe",x"87",x"c8"),
   192 => (x"c1",x"48",x"c0",x"87"),
   193 => (x"da",x"fa",x"87",x"e2"),
   194 => (x"cf",x"49",x"70",x"87"),
   195 => (x"c6",x"99",x"ff",x"ff"),
   196 => (x"c8",x"02",x"a9",x"ea"),
   197 => (x"87",x"d3",x"fe",x"87"),
   198 => (x"cb",x"c1",x"48",x"c0"),
   199 => (x"7c",x"ff",x"c3",x"87"),
   200 => (x"fc",x"4b",x"f1",x"c0"),
   201 => (x"98",x"70",x"87",x"f4"),
   202 => (x"87",x"eb",x"c0",x"02"),
   203 => (x"ff",x"c0",x"1e",x"c0"),
   204 => (x"49",x"fa",x"c1",x"f0"),
   205 => (x"c4",x"87",x"de",x"fa"),
   206 => (x"05",x"98",x"70",x"86"),
   207 => (x"ff",x"c3",x"87",x"d9"),
   208 => (x"c3",x"49",x"6c",x"7c"),
   209 => (x"7c",x"7c",x"7c",x"ff"),
   210 => (x"99",x"c0",x"c1",x"7c"),
   211 => (x"c1",x"87",x"c4",x"02"),
   212 => (x"c0",x"87",x"d5",x"48"),
   213 => (x"c2",x"87",x"d1",x"48"),
   214 => (x"87",x"c4",x"05",x"ab"),
   215 => (x"87",x"c8",x"48",x"c0"),
   216 => (x"fe",x"05",x"8b",x"c1"),
   217 => (x"48",x"c0",x"87",x"fd"),
   218 => (x"1e",x"87",x"e4",x"f9"),
   219 => (x"ef",x"c3",x"1e",x"73"),
   220 => (x"78",x"c1",x"48",x"ec"),
   221 => (x"d0",x"ff",x"4b",x"c7"),
   222 => (x"fb",x"78",x"c2",x"48"),
   223 => (x"d0",x"ff",x"87",x"c8"),
   224 => (x"c0",x"78",x"c3",x"48"),
   225 => (x"d0",x"e5",x"c0",x"1e"),
   226 => (x"f9",x"49",x"c0",x"c1"),
   227 => (x"86",x"c4",x"87",x"c7"),
   228 => (x"c1",x"05",x"a8",x"c1"),
   229 => (x"ab",x"c2",x"4b",x"87"),
   230 => (x"c0",x"87",x"c5",x"05"),
   231 => (x"87",x"f9",x"c0",x"48"),
   232 => (x"ff",x"05",x"8b",x"c1"),
   233 => (x"f7",x"fc",x"87",x"d0"),
   234 => (x"f0",x"ef",x"c3",x"87"),
   235 => (x"05",x"98",x"70",x"58"),
   236 => (x"1e",x"c1",x"87",x"cd"),
   237 => (x"c1",x"f0",x"ff",x"c0"),
   238 => (x"d8",x"f8",x"49",x"d0"),
   239 => (x"ff",x"86",x"c4",x"87"),
   240 => (x"ff",x"c3",x"48",x"d4"),
   241 => (x"87",x"e0",x"c4",x"78"),
   242 => (x"58",x"f4",x"ef",x"c3"),
   243 => (x"c2",x"48",x"d0",x"ff"),
   244 => (x"48",x"d4",x"ff",x"78"),
   245 => (x"c1",x"78",x"ff",x"c3"),
   246 => (x"87",x"f5",x"f7",x"48"),
   247 => (x"5c",x"5b",x"5e",x"0e"),
   248 => (x"4a",x"71",x"0e",x"5d"),
   249 => (x"ff",x"4d",x"ff",x"c3"),
   250 => (x"7c",x"75",x"4c",x"d4"),
   251 => (x"c4",x"48",x"d0",x"ff"),
   252 => (x"7c",x"75",x"78",x"c3"),
   253 => (x"ff",x"c0",x"1e",x"72"),
   254 => (x"49",x"d8",x"c1",x"f0"),
   255 => (x"c4",x"87",x"d6",x"f7"),
   256 => (x"02",x"98",x"70",x"86"),
   257 => (x"48",x"c0",x"87",x"c5"),
   258 => (x"75",x"87",x"f0",x"c0"),
   259 => (x"7c",x"fe",x"c3",x"7c"),
   260 => (x"d4",x"1e",x"c0",x"c8"),
   261 => (x"dc",x"f5",x"49",x"66"),
   262 => (x"75",x"86",x"c4",x"87"),
   263 => (x"75",x"7c",x"75",x"7c"),
   264 => (x"e0",x"da",x"d8",x"7c"),
   265 => (x"6c",x"7c",x"75",x"4b"),
   266 => (x"c5",x"05",x"99",x"49"),
   267 => (x"05",x"8b",x"c1",x"87"),
   268 => (x"7c",x"75",x"87",x"f3"),
   269 => (x"c2",x"48",x"d0",x"ff"),
   270 => (x"f6",x"48",x"c1",x"78"),
   271 => (x"ff",x"1e",x"87",x"cf"),
   272 => (x"d0",x"ff",x"4a",x"d4"),
   273 => (x"78",x"d1",x"c4",x"48"),
   274 => (x"c1",x"7a",x"ff",x"c3"),
   275 => (x"87",x"f8",x"05",x"89"),
   276 => (x"73",x"1e",x"4f",x"26"),
   277 => (x"c5",x"4b",x"71",x"1e"),
   278 => (x"4a",x"df",x"cd",x"ee"),
   279 => (x"c3",x"48",x"d4",x"ff"),
   280 => (x"48",x"68",x"78",x"ff"),
   281 => (x"02",x"a8",x"fe",x"c3"),
   282 => (x"8a",x"c1",x"87",x"c5"),
   283 => (x"72",x"87",x"ed",x"05"),
   284 => (x"87",x"c5",x"05",x"9a"),
   285 => (x"ea",x"c0",x"48",x"c0"),
   286 => (x"02",x"9b",x"73",x"87"),
   287 => (x"66",x"c8",x"87",x"cc"),
   288 => (x"f4",x"49",x"73",x"1e"),
   289 => (x"86",x"c4",x"87",x"c5"),
   290 => (x"66",x"c8",x"87",x"c6"),
   291 => (x"87",x"ee",x"fe",x"49"),
   292 => (x"c3",x"48",x"d4",x"ff"),
   293 => (x"73",x"78",x"78",x"ff"),
   294 => (x"87",x"c5",x"05",x"9b"),
   295 => (x"d0",x"48",x"d0",x"ff"),
   296 => (x"f4",x"48",x"c1",x"78"),
   297 => (x"73",x"1e",x"87",x"eb"),
   298 => (x"c0",x"4a",x"71",x"1e"),
   299 => (x"48",x"d4",x"ff",x"4b"),
   300 => (x"ff",x"78",x"ff",x"c3"),
   301 => (x"c3",x"c4",x"48",x"d0"),
   302 => (x"48",x"d4",x"ff",x"78"),
   303 => (x"72",x"78",x"ff",x"c3"),
   304 => (x"f0",x"ff",x"c0",x"1e"),
   305 => (x"f4",x"49",x"d1",x"c1"),
   306 => (x"86",x"c4",x"87",x"cb"),
   307 => (x"cd",x"05",x"98",x"70"),
   308 => (x"1e",x"c0",x"c8",x"87"),
   309 => (x"fd",x"49",x"66",x"cc"),
   310 => (x"86",x"c4",x"87",x"f8"),
   311 => (x"d0",x"ff",x"4b",x"70"),
   312 => (x"73",x"78",x"c2",x"48"),
   313 => (x"87",x"e9",x"f3",x"48"),
   314 => (x"5c",x"5b",x"5e",x"0e"),
   315 => (x"1e",x"c0",x"0e",x"5d"),
   316 => (x"c1",x"f0",x"ff",x"c0"),
   317 => (x"dc",x"f3",x"49",x"c9"),
   318 => (x"c3",x"1e",x"d2",x"87"),
   319 => (x"fd",x"49",x"f4",x"ef"),
   320 => (x"86",x"c8",x"87",x"d0"),
   321 => (x"84",x"c1",x"4c",x"c0"),
   322 => (x"04",x"ac",x"b7",x"d2"),
   323 => (x"ef",x"c3",x"87",x"f8"),
   324 => (x"49",x"bf",x"97",x"f4"),
   325 => (x"c1",x"99",x"c0",x"c3"),
   326 => (x"c0",x"05",x"a9",x"c0"),
   327 => (x"ef",x"c3",x"87",x"e7"),
   328 => (x"49",x"bf",x"97",x"fb"),
   329 => (x"ef",x"c3",x"31",x"d0"),
   330 => (x"4a",x"bf",x"97",x"fc"),
   331 => (x"b1",x"72",x"32",x"c8"),
   332 => (x"97",x"fd",x"ef",x"c3"),
   333 => (x"71",x"b1",x"4a",x"bf"),
   334 => (x"ff",x"ff",x"cf",x"4c"),
   335 => (x"84",x"c1",x"9c",x"ff"),
   336 => (x"e7",x"c1",x"34",x"ca"),
   337 => (x"fd",x"ef",x"c3",x"87"),
   338 => (x"c1",x"49",x"bf",x"97"),
   339 => (x"c3",x"99",x"c6",x"31"),
   340 => (x"bf",x"97",x"fe",x"ef"),
   341 => (x"2a",x"b7",x"c7",x"4a"),
   342 => (x"ef",x"c3",x"b1",x"72"),
   343 => (x"4a",x"bf",x"97",x"f9"),
   344 => (x"c3",x"9d",x"cf",x"4d"),
   345 => (x"bf",x"97",x"fa",x"ef"),
   346 => (x"ca",x"9a",x"c3",x"4a"),
   347 => (x"fb",x"ef",x"c3",x"32"),
   348 => (x"c2",x"4b",x"bf",x"97"),
   349 => (x"c3",x"b2",x"73",x"33"),
   350 => (x"bf",x"97",x"fc",x"ef"),
   351 => (x"9b",x"c0",x"c3",x"4b"),
   352 => (x"73",x"2b",x"b7",x"c6"),
   353 => (x"c1",x"81",x"c2",x"b2"),
   354 => (x"70",x"30",x"71",x"48"),
   355 => (x"75",x"48",x"c1",x"49"),
   356 => (x"72",x"4d",x"70",x"30"),
   357 => (x"71",x"84",x"c1",x"4c"),
   358 => (x"b7",x"c0",x"c8",x"94"),
   359 => (x"87",x"cc",x"06",x"ad"),
   360 => (x"2d",x"b7",x"34",x"c1"),
   361 => (x"ad",x"b7",x"c0",x"c8"),
   362 => (x"87",x"f4",x"ff",x"01"),
   363 => (x"dc",x"f0",x"48",x"74"),
   364 => (x"5b",x"5e",x"0e",x"87"),
   365 => (x"f8",x"0e",x"5d",x"5c"),
   366 => (x"da",x"f8",x"c3",x"86"),
   367 => (x"c3",x"78",x"c0",x"48"),
   368 => (x"c0",x"1e",x"d2",x"f0"),
   369 => (x"87",x"de",x"fb",x"49"),
   370 => (x"98",x"70",x"86",x"c4"),
   371 => (x"c0",x"87",x"c5",x"05"),
   372 => (x"87",x"ce",x"c9",x"48"),
   373 => (x"7e",x"c1",x"4d",x"c0"),
   374 => (x"bf",x"f0",x"fb",x"c0"),
   375 => (x"c8",x"f1",x"c3",x"49"),
   376 => (x"4b",x"c8",x"71",x"4a"),
   377 => (x"70",x"87",x"c1",x"eb"),
   378 => (x"87",x"c2",x"05",x"98"),
   379 => (x"fb",x"c0",x"7e",x"c0"),
   380 => (x"c3",x"49",x"bf",x"ec"),
   381 => (x"71",x"4a",x"e4",x"f1"),
   382 => (x"eb",x"ea",x"4b",x"c8"),
   383 => (x"05",x"98",x"70",x"87"),
   384 => (x"7e",x"c0",x"87",x"c2"),
   385 => (x"fd",x"c0",x"02",x"6e"),
   386 => (x"d8",x"f7",x"c3",x"87"),
   387 => (x"f8",x"c3",x"4d",x"bf"),
   388 => (x"7e",x"bf",x"9f",x"d0"),
   389 => (x"ea",x"d6",x"c5",x"48"),
   390 => (x"87",x"c7",x"05",x"a8"),
   391 => (x"bf",x"d8",x"f7",x"c3"),
   392 => (x"6e",x"87",x"ce",x"4d"),
   393 => (x"d5",x"e9",x"ca",x"48"),
   394 => (x"87",x"c5",x"02",x"a8"),
   395 => (x"f1",x"c7",x"48",x"c0"),
   396 => (x"d2",x"f0",x"c3",x"87"),
   397 => (x"f9",x"49",x"75",x"1e"),
   398 => (x"86",x"c4",x"87",x"ec"),
   399 => (x"c5",x"05",x"98",x"70"),
   400 => (x"c7",x"48",x"c0",x"87"),
   401 => (x"fb",x"c0",x"87",x"dc"),
   402 => (x"c3",x"49",x"bf",x"ec"),
   403 => (x"71",x"4a",x"e4",x"f1"),
   404 => (x"d3",x"e9",x"4b",x"c8"),
   405 => (x"05",x"98",x"70",x"87"),
   406 => (x"f8",x"c3",x"87",x"c8"),
   407 => (x"78",x"c1",x"48",x"da"),
   408 => (x"fb",x"c0",x"87",x"da"),
   409 => (x"c3",x"49",x"bf",x"f0"),
   410 => (x"71",x"4a",x"c8",x"f1"),
   411 => (x"f7",x"e8",x"4b",x"c8"),
   412 => (x"02",x"98",x"70",x"87"),
   413 => (x"c0",x"87",x"c5",x"c0"),
   414 => (x"87",x"e6",x"c6",x"48"),
   415 => (x"97",x"d0",x"f8",x"c3"),
   416 => (x"d5",x"c1",x"49",x"bf"),
   417 => (x"cd",x"c0",x"05",x"a9"),
   418 => (x"d1",x"f8",x"c3",x"87"),
   419 => (x"c2",x"49",x"bf",x"97"),
   420 => (x"c0",x"02",x"a9",x"ea"),
   421 => (x"48",x"c0",x"87",x"c5"),
   422 => (x"c3",x"87",x"c7",x"c6"),
   423 => (x"bf",x"97",x"d2",x"f0"),
   424 => (x"e9",x"c3",x"48",x"7e"),
   425 => (x"ce",x"c0",x"02",x"a8"),
   426 => (x"c3",x"48",x"6e",x"87"),
   427 => (x"c0",x"02",x"a8",x"eb"),
   428 => (x"48",x"c0",x"87",x"c5"),
   429 => (x"c3",x"87",x"eb",x"c5"),
   430 => (x"bf",x"97",x"dd",x"f0"),
   431 => (x"c0",x"05",x"99",x"49"),
   432 => (x"f0",x"c3",x"87",x"cc"),
   433 => (x"49",x"bf",x"97",x"de"),
   434 => (x"c0",x"02",x"a9",x"c2"),
   435 => (x"48",x"c0",x"87",x"c5"),
   436 => (x"c3",x"87",x"cf",x"c5"),
   437 => (x"bf",x"97",x"df",x"f0"),
   438 => (x"d6",x"f8",x"c3",x"48"),
   439 => (x"48",x"4c",x"70",x"58"),
   440 => (x"f8",x"c3",x"88",x"c1"),
   441 => (x"f0",x"c3",x"58",x"da"),
   442 => (x"49",x"bf",x"97",x"e0"),
   443 => (x"f0",x"c3",x"81",x"75"),
   444 => (x"4a",x"bf",x"97",x"e1"),
   445 => (x"a1",x"72",x"32",x"c8"),
   446 => (x"e7",x"fc",x"c3",x"7e"),
   447 => (x"c3",x"78",x"6e",x"48"),
   448 => (x"bf",x"97",x"e2",x"f0"),
   449 => (x"58",x"a6",x"c8",x"48"),
   450 => (x"bf",x"da",x"f8",x"c3"),
   451 => (x"87",x"d4",x"c2",x"02"),
   452 => (x"bf",x"ec",x"fb",x"c0"),
   453 => (x"e4",x"f1",x"c3",x"49"),
   454 => (x"4b",x"c8",x"71",x"4a"),
   455 => (x"70",x"87",x"c9",x"e6"),
   456 => (x"c5",x"c0",x"02",x"98"),
   457 => (x"c3",x"48",x"c0",x"87"),
   458 => (x"f8",x"c3",x"87",x"f8"),
   459 => (x"c3",x"4c",x"bf",x"d2"),
   460 => (x"c3",x"5c",x"fb",x"fc"),
   461 => (x"bf",x"97",x"f7",x"f0"),
   462 => (x"c3",x"31",x"c8",x"49"),
   463 => (x"bf",x"97",x"f6",x"f0"),
   464 => (x"c3",x"49",x"a1",x"4a"),
   465 => (x"bf",x"97",x"f8",x"f0"),
   466 => (x"72",x"32",x"d0",x"4a"),
   467 => (x"f0",x"c3",x"49",x"a1"),
   468 => (x"4a",x"bf",x"97",x"f9"),
   469 => (x"a1",x"72",x"32",x"d8"),
   470 => (x"91",x"66",x"c4",x"49"),
   471 => (x"bf",x"e7",x"fc",x"c3"),
   472 => (x"ef",x"fc",x"c3",x"81"),
   473 => (x"ff",x"f0",x"c3",x"59"),
   474 => (x"c8",x"4a",x"bf",x"97"),
   475 => (x"fe",x"f0",x"c3",x"32"),
   476 => (x"a2",x"4b",x"bf",x"97"),
   477 => (x"c0",x"f1",x"c3",x"4a"),
   478 => (x"d0",x"4b",x"bf",x"97"),
   479 => (x"4a",x"a2",x"73",x"33"),
   480 => (x"97",x"c1",x"f1",x"c3"),
   481 => (x"9b",x"cf",x"4b",x"bf"),
   482 => (x"a2",x"73",x"33",x"d8"),
   483 => (x"f3",x"fc",x"c3",x"4a"),
   484 => (x"ef",x"fc",x"c3",x"5a"),
   485 => (x"8a",x"c2",x"4a",x"bf"),
   486 => (x"fc",x"c3",x"92",x"74"),
   487 => (x"a1",x"72",x"48",x"f3"),
   488 => (x"87",x"ca",x"c1",x"78"),
   489 => (x"97",x"e4",x"f0",x"c3"),
   490 => (x"31",x"c8",x"49",x"bf"),
   491 => (x"97",x"e3",x"f0",x"c3"),
   492 => (x"49",x"a1",x"4a",x"bf"),
   493 => (x"59",x"e2",x"f8",x"c3"),
   494 => (x"bf",x"de",x"f8",x"c3"),
   495 => (x"c7",x"31",x"c5",x"49"),
   496 => (x"29",x"c9",x"81",x"ff"),
   497 => (x"59",x"fb",x"fc",x"c3"),
   498 => (x"97",x"e9",x"f0",x"c3"),
   499 => (x"32",x"c8",x"4a",x"bf"),
   500 => (x"97",x"e8",x"f0",x"c3"),
   501 => (x"4a",x"a2",x"4b",x"bf"),
   502 => (x"6e",x"92",x"66",x"c4"),
   503 => (x"f7",x"fc",x"c3",x"82"),
   504 => (x"ef",x"fc",x"c3",x"5a"),
   505 => (x"c3",x"78",x"c0",x"48"),
   506 => (x"72",x"48",x"eb",x"fc"),
   507 => (x"fc",x"c3",x"78",x"a1"),
   508 => (x"fc",x"c3",x"48",x"fb"),
   509 => (x"c3",x"78",x"bf",x"ef"),
   510 => (x"c3",x"48",x"ff",x"fc"),
   511 => (x"78",x"bf",x"f3",x"fc"),
   512 => (x"bf",x"da",x"f8",x"c3"),
   513 => (x"87",x"c9",x"c0",x"02"),
   514 => (x"30",x"c4",x"48",x"74"),
   515 => (x"c9",x"c0",x"7e",x"70"),
   516 => (x"f7",x"fc",x"c3",x"87"),
   517 => (x"30",x"c4",x"48",x"bf"),
   518 => (x"f8",x"c3",x"7e",x"70"),
   519 => (x"78",x"6e",x"48",x"de"),
   520 => (x"8e",x"f8",x"48",x"c1"),
   521 => (x"4c",x"26",x"4d",x"26"),
   522 => (x"4f",x"26",x"4b",x"26"),
   523 => (x"5c",x"5b",x"5e",x"0e"),
   524 => (x"4a",x"71",x"0e",x"5d"),
   525 => (x"bf",x"da",x"f8",x"c3"),
   526 => (x"72",x"87",x"cb",x"02"),
   527 => (x"72",x"2b",x"c7",x"4b"),
   528 => (x"9c",x"ff",x"c1",x"4c"),
   529 => (x"4b",x"72",x"87",x"c9"),
   530 => (x"4c",x"72",x"2b",x"c8"),
   531 => (x"c3",x"9c",x"ff",x"c3"),
   532 => (x"83",x"bf",x"e7",x"fc"),
   533 => (x"bf",x"e8",x"fb",x"c0"),
   534 => (x"87",x"d9",x"02",x"ab"),
   535 => (x"5b",x"ec",x"fb",x"c0"),
   536 => (x"1e",x"d2",x"f0",x"c3"),
   537 => (x"fd",x"f0",x"49",x"73"),
   538 => (x"70",x"86",x"c4",x"87"),
   539 => (x"87",x"c5",x"05",x"98"),
   540 => (x"e6",x"c0",x"48",x"c0"),
   541 => (x"da",x"f8",x"c3",x"87"),
   542 => (x"87",x"d2",x"02",x"bf"),
   543 => (x"91",x"c4",x"49",x"74"),
   544 => (x"81",x"d2",x"f0",x"c3"),
   545 => (x"ff",x"cf",x"4d",x"69"),
   546 => (x"9d",x"ff",x"ff",x"ff"),
   547 => (x"49",x"74",x"87",x"cb"),
   548 => (x"f0",x"c3",x"91",x"c2"),
   549 => (x"69",x"9f",x"81",x"d2"),
   550 => (x"fe",x"48",x"75",x"4d"),
   551 => (x"5e",x"0e",x"87",x"c6"),
   552 => (x"0e",x"5d",x"5c",x"5b"),
   553 => (x"c0",x"4d",x"71",x"1e"),
   554 => (x"d1",x"49",x"c1",x"1e"),
   555 => (x"86",x"c4",x"87",x"e2"),
   556 => (x"02",x"9c",x"4c",x"70"),
   557 => (x"c3",x"87",x"c2",x"c1"),
   558 => (x"75",x"4a",x"e2",x"f8"),
   559 => (x"cc",x"df",x"ff",x"49"),
   560 => (x"02",x"98",x"70",x"87"),
   561 => (x"74",x"87",x"f2",x"c0"),
   562 => (x"cb",x"49",x"75",x"4a"),
   563 => (x"f1",x"df",x"ff",x"4b"),
   564 => (x"02",x"98",x"70",x"87"),
   565 => (x"c0",x"87",x"e2",x"c0"),
   566 => (x"02",x"9c",x"74",x"1e"),
   567 => (x"a6",x"c4",x"87",x"c7"),
   568 => (x"c5",x"78",x"c0",x"48"),
   569 => (x"48",x"a6",x"c4",x"87"),
   570 => (x"66",x"c4",x"78",x"c1"),
   571 => (x"87",x"e0",x"d0",x"49"),
   572 => (x"4c",x"70",x"86",x"c4"),
   573 => (x"fe",x"fe",x"05",x"9c"),
   574 => (x"26",x"48",x"74",x"87"),
   575 => (x"0e",x"87",x"e5",x"fc"),
   576 => (x"5d",x"5c",x"5b",x"5e"),
   577 => (x"71",x"86",x"f8",x"0e"),
   578 => (x"c5",x"05",x"9b",x"4b"),
   579 => (x"c2",x"48",x"c0",x"87"),
   580 => (x"a3",x"c8",x"87",x"d4"),
   581 => (x"d8",x"7d",x"c0",x"4d"),
   582 => (x"87",x"c7",x"02",x"66"),
   583 => (x"bf",x"97",x"66",x"d8"),
   584 => (x"c0",x"87",x"c5",x"05"),
   585 => (x"87",x"fe",x"c1",x"48"),
   586 => (x"fd",x"49",x"66",x"d8"),
   587 => (x"7e",x"70",x"87",x"f0"),
   588 => (x"ef",x"c1",x"02",x"6e"),
   589 => (x"dc",x"49",x"6e",x"87"),
   590 => (x"6e",x"7d",x"69",x"81"),
   591 => (x"c4",x"81",x"da",x"49"),
   592 => (x"69",x"9f",x"4c",x"a3"),
   593 => (x"da",x"f8",x"c3",x"7c"),
   594 => (x"87",x"d0",x"02",x"bf"),
   595 => (x"81",x"d4",x"49",x"6e"),
   596 => (x"4a",x"49",x"69",x"9f"),
   597 => (x"9a",x"ff",x"ff",x"c0"),
   598 => (x"87",x"c2",x"32",x"d0"),
   599 => (x"49",x"72",x"4a",x"c0"),
   600 => (x"70",x"80",x"6c",x"48"),
   601 => (x"cc",x"7b",x"c0",x"7c"),
   602 => (x"79",x"6c",x"49",x"a3"),
   603 => (x"c0",x"49",x"a3",x"d0"),
   604 => (x"48",x"a6",x"c4",x"79"),
   605 => (x"a3",x"d4",x"78",x"c0"),
   606 => (x"49",x"66",x"c4",x"4a"),
   607 => (x"a1",x"72",x"91",x"c8"),
   608 => (x"6c",x"41",x"c0",x"49"),
   609 => (x"48",x"66",x"c4",x"79"),
   610 => (x"a6",x"c8",x"80",x"c1"),
   611 => (x"a8",x"b7",x"d0",x"58"),
   612 => (x"87",x"e2",x"ff",x"04"),
   613 => (x"2a",x"c9",x"4a",x"6d"),
   614 => (x"d4",x"c2",x"2a",x"c7"),
   615 => (x"79",x"72",x"49",x"a3"),
   616 => (x"87",x"c2",x"48",x"6e"),
   617 => (x"8e",x"f8",x"48",x"c0"),
   618 => (x"0e",x"87",x"f9",x"f9"),
   619 => (x"5d",x"5c",x"5b",x"5e"),
   620 => (x"c0",x"4c",x"71",x"0e"),
   621 => (x"ff",x"48",x"e8",x"fb"),
   622 => (x"02",x"9c",x"74",x"78"),
   623 => (x"c8",x"87",x"ca",x"c1"),
   624 => (x"02",x"69",x"49",x"a4"),
   625 => (x"d0",x"87",x"c2",x"c1"),
   626 => (x"49",x"6c",x"4a",x"66"),
   627 => (x"5a",x"a6",x"d4",x"82"),
   628 => (x"b9",x"4d",x"66",x"d0"),
   629 => (x"bf",x"d6",x"f8",x"c3"),
   630 => (x"72",x"ba",x"ff",x"4a"),
   631 => (x"02",x"99",x"71",x"99"),
   632 => (x"c4",x"87",x"e4",x"c0"),
   633 => (x"49",x"6b",x"4b",x"a4"),
   634 => (x"70",x"87",x"c1",x"f9"),
   635 => (x"d2",x"f8",x"c3",x"7b"),
   636 => (x"81",x"6c",x"49",x"bf"),
   637 => (x"b9",x"75",x"7c",x"71"),
   638 => (x"bf",x"d6",x"f8",x"c3"),
   639 => (x"72",x"ba",x"ff",x"4a"),
   640 => (x"05",x"99",x"71",x"99"),
   641 => (x"75",x"87",x"dc",x"ff"),
   642 => (x"87",x"d8",x"f8",x"7c"),
   643 => (x"71",x"1e",x"73",x"1e"),
   644 => (x"c7",x"02",x"9b",x"4b"),
   645 => (x"49",x"a3",x"c8",x"87"),
   646 => (x"87",x"c5",x"05",x"69"),
   647 => (x"eb",x"c0",x"48",x"c0"),
   648 => (x"eb",x"fc",x"c3",x"87"),
   649 => (x"a3",x"c4",x"4a",x"bf"),
   650 => (x"c2",x"49",x"69",x"49"),
   651 => (x"d2",x"f8",x"c3",x"89"),
   652 => (x"a2",x"71",x"91",x"bf"),
   653 => (x"d6",x"f8",x"c3",x"4a"),
   654 => (x"99",x"6b",x"49",x"bf"),
   655 => (x"c8",x"4a",x"a2",x"71"),
   656 => (x"49",x"72",x"1e",x"66"),
   657 => (x"c4",x"87",x"df",x"e9"),
   658 => (x"48",x"49",x"70",x"86"),
   659 => (x"1e",x"87",x"d9",x"f7"),
   660 => (x"4b",x"71",x"1e",x"73"),
   661 => (x"87",x"c7",x"02",x"9b"),
   662 => (x"69",x"49",x"a3",x"c8"),
   663 => (x"c0",x"87",x"c5",x"05"),
   664 => (x"87",x"eb",x"c0",x"48"),
   665 => (x"bf",x"eb",x"fc",x"c3"),
   666 => (x"49",x"a3",x"c4",x"4a"),
   667 => (x"89",x"c2",x"49",x"69"),
   668 => (x"bf",x"d2",x"f8",x"c3"),
   669 => (x"4a",x"a2",x"71",x"91"),
   670 => (x"bf",x"d6",x"f8",x"c3"),
   671 => (x"71",x"99",x"6b",x"49"),
   672 => (x"66",x"c8",x"4a",x"a2"),
   673 => (x"e5",x"49",x"72",x"1e"),
   674 => (x"86",x"c4",x"87",x"d2"),
   675 => (x"f6",x"48",x"49",x"70"),
   676 => (x"5e",x"0e",x"87",x"d6"),
   677 => (x"0e",x"5d",x"5c",x"5b"),
   678 => (x"4b",x"71",x"86",x"f8"),
   679 => (x"ff",x"48",x"a6",x"c4"),
   680 => (x"49",x"a3",x"c8",x"78"),
   681 => (x"4c",x"c0",x"4d",x"69"),
   682 => (x"74",x"4a",x"a3",x"d4"),
   683 => (x"72",x"91",x"c8",x"49"),
   684 => (x"49",x"69",x"49",x"a1"),
   685 => (x"71",x"48",x"66",x"d8"),
   686 => (x"d8",x"7e",x"70",x"88"),
   687 => (x"ca",x"01",x"a9",x"66"),
   688 => (x"06",x"ad",x"6e",x"87"),
   689 => (x"a6",x"c8",x"87",x"c5"),
   690 => (x"c1",x"4d",x"6e",x"5c"),
   691 => (x"ac",x"b7",x"d0",x"84"),
   692 => (x"87",x"d4",x"ff",x"04"),
   693 => (x"f8",x"48",x"66",x"c4"),
   694 => (x"87",x"c8",x"f5",x"8e"),
   695 => (x"5c",x"5b",x"5e",x"0e"),
   696 => (x"86",x"ec",x"0e",x"5d"),
   697 => (x"c8",x"59",x"a6",x"c8"),
   698 => (x"ff",x"c1",x"48",x"a6"),
   699 => (x"ff",x"ff",x"ff",x"ff"),
   700 => (x"ff",x"80",x"c4",x"78"),
   701 => (x"c0",x"4d",x"c0",x"78"),
   702 => (x"4b",x"66",x"c4",x"4c"),
   703 => (x"49",x"74",x"83",x"d4"),
   704 => (x"a1",x"73",x"91",x"c8"),
   705 => (x"c8",x"4a",x"75",x"49"),
   706 => (x"7e",x"a2",x"73",x"92"),
   707 => (x"bf",x"6e",x"49",x"69"),
   708 => (x"59",x"a6",x"d4",x"89"),
   709 => (x"c6",x"05",x"ad",x"74"),
   710 => (x"48",x"a6",x"d0",x"87"),
   711 => (x"d0",x"78",x"bf",x"6e"),
   712 => (x"b7",x"c0",x"48",x"66"),
   713 => (x"87",x"cf",x"04",x"a8"),
   714 => (x"c8",x"49",x"66",x"d0"),
   715 => (x"c6",x"03",x"a9",x"66"),
   716 => (x"5c",x"a6",x"d0",x"87"),
   717 => (x"c1",x"59",x"a6",x"cc"),
   718 => (x"ac",x"b7",x"d0",x"84"),
   719 => (x"87",x"f9",x"fe",x"04"),
   720 => (x"b7",x"d0",x"85",x"c1"),
   721 => (x"ee",x"fe",x"04",x"ad"),
   722 => (x"48",x"66",x"cc",x"87"),
   723 => (x"d3",x"f3",x"8e",x"ec"),
   724 => (x"5b",x"5e",x"0e",x"87"),
   725 => (x"4b",x"71",x"0e",x"5c"),
   726 => (x"a3",x"c8",x"4c",x"c0"),
   727 => (x"c4",x"49",x"69",x"49"),
   728 => (x"91",x"4a",x"74",x"29"),
   729 => (x"49",x"73",x"1e",x"71"),
   730 => (x"86",x"c4",x"87",x"d4"),
   731 => (x"b7",x"d0",x"84",x"c1"),
   732 => (x"87",x"e6",x"04",x"ac"),
   733 => (x"49",x"73",x"1e",x"c0"),
   734 => (x"f2",x"26",x"87",x"c4"),
   735 => (x"5e",x"0e",x"87",x"e8"),
   736 => (x"0e",x"5d",x"5c",x"5b"),
   737 => (x"4b",x"71",x"86",x"f0"),
   738 => (x"4c",x"66",x"e0",x"c0"),
   739 => (x"9b",x"73",x"2c",x"c9"),
   740 => (x"87",x"e1",x"c3",x"02"),
   741 => (x"69",x"49",x"a3",x"c8"),
   742 => (x"87",x"d9",x"c3",x"02"),
   743 => (x"c0",x"49",x"a3",x"d0"),
   744 => (x"6b",x"79",x"66",x"e0"),
   745 => (x"c3",x"02",x"ac",x"7e"),
   746 => (x"f8",x"c3",x"87",x"cb"),
   747 => (x"ff",x"49",x"bf",x"d6"),
   748 => (x"74",x"4a",x"71",x"b9"),
   749 => (x"6e",x"48",x"71",x"9a"),
   750 => (x"58",x"a6",x"cc",x"98"),
   751 => (x"c4",x"4d",x"a3",x"c4"),
   752 => (x"78",x"6d",x"48",x"a6"),
   753 => (x"05",x"aa",x"66",x"c8"),
   754 => (x"7b",x"74",x"87",x"c5"),
   755 => (x"72",x"87",x"d1",x"c2"),
   756 => (x"fa",x"49",x"73",x"1e"),
   757 => (x"86",x"c4",x"87",x"fc"),
   758 => (x"c0",x"48",x"7e",x"70"),
   759 => (x"d0",x"04",x"a8",x"b7"),
   760 => (x"4a",x"a3",x"d4",x"87"),
   761 => (x"91",x"c8",x"49",x"6e"),
   762 => (x"21",x"49",x"a1",x"72"),
   763 => (x"c7",x"7d",x"69",x"7b"),
   764 => (x"cc",x"7b",x"c0",x"87"),
   765 => (x"7d",x"69",x"49",x"a3"),
   766 => (x"73",x"1e",x"66",x"c8"),
   767 => (x"87",x"d2",x"fa",x"49"),
   768 => (x"7e",x"70",x"86",x"c4"),
   769 => (x"49",x"a3",x"d4",x"c2"),
   770 => (x"69",x"48",x"a6",x"cc"),
   771 => (x"48",x"66",x"c8",x"78"),
   772 => (x"06",x"a8",x"66",x"cc"),
   773 => (x"48",x"6e",x"87",x"c9"),
   774 => (x"04",x"a8",x"b7",x"c0"),
   775 => (x"6e",x"87",x"e0",x"c0"),
   776 => (x"a8",x"b7",x"c0",x"48"),
   777 => (x"87",x"ec",x"c0",x"04"),
   778 => (x"6e",x"4a",x"a3",x"d4"),
   779 => (x"72",x"91",x"c8",x"49"),
   780 => (x"66",x"c8",x"49",x"a1"),
   781 => (x"70",x"88",x"69",x"48"),
   782 => (x"a9",x"66",x"cc",x"49"),
   783 => (x"73",x"87",x"d5",x"06"),
   784 => (x"87",x"d8",x"fa",x"49"),
   785 => (x"a3",x"d4",x"49",x"70"),
   786 => (x"72",x"91",x"c8",x"4a"),
   787 => (x"66",x"c8",x"49",x"a1"),
   788 => (x"79",x"66",x"c4",x"41"),
   789 => (x"49",x"74",x"8c",x"6b"),
   790 => (x"f5",x"49",x"73",x"1e"),
   791 => (x"86",x"c4",x"87",x"cd"),
   792 => (x"49",x"66",x"e0",x"c0"),
   793 => (x"02",x"99",x"ff",x"c7"),
   794 => (x"f0",x"c3",x"87",x"cb"),
   795 => (x"49",x"73",x"1e",x"d2"),
   796 => (x"c4",x"87",x"d9",x"f6"),
   797 => (x"ee",x"8e",x"f0",x"86"),
   798 => (x"73",x"1e",x"87",x"ea"),
   799 => (x"9b",x"4b",x"71",x"1e"),
   800 => (x"87",x"e4",x"c0",x"02"),
   801 => (x"5b",x"ff",x"fc",x"c3"),
   802 => (x"8a",x"c2",x"4a",x"73"),
   803 => (x"bf",x"d2",x"f8",x"c3"),
   804 => (x"fc",x"c3",x"92",x"49"),
   805 => (x"72",x"48",x"bf",x"eb"),
   806 => (x"c3",x"fd",x"c3",x"80"),
   807 => (x"c4",x"48",x"71",x"58"),
   808 => (x"e2",x"f8",x"c3",x"30"),
   809 => (x"87",x"ed",x"c0",x"58"),
   810 => (x"48",x"fb",x"fc",x"c3"),
   811 => (x"bf",x"ef",x"fc",x"c3"),
   812 => (x"ff",x"fc",x"c3",x"78"),
   813 => (x"f3",x"fc",x"c3",x"48"),
   814 => (x"f8",x"c3",x"78",x"bf"),
   815 => (x"c9",x"02",x"bf",x"da"),
   816 => (x"d2",x"f8",x"c3",x"87"),
   817 => (x"31",x"c4",x"49",x"bf"),
   818 => (x"fc",x"c3",x"87",x"c7"),
   819 => (x"c4",x"49",x"bf",x"f7"),
   820 => (x"e2",x"f8",x"c3",x"31"),
   821 => (x"87",x"d0",x"ed",x"59"),
   822 => (x"5c",x"5b",x"5e",x"0e"),
   823 => (x"c0",x"4a",x"71",x"0e"),
   824 => (x"02",x"9a",x"72",x"4b"),
   825 => (x"da",x"87",x"e1",x"c0"),
   826 => (x"69",x"9f",x"49",x"a2"),
   827 => (x"da",x"f8",x"c3",x"4b"),
   828 => (x"87",x"cf",x"02",x"bf"),
   829 => (x"9f",x"49",x"a2",x"d4"),
   830 => (x"c0",x"4c",x"49",x"69"),
   831 => (x"d0",x"9c",x"ff",x"ff"),
   832 => (x"c0",x"87",x"c2",x"34"),
   833 => (x"b3",x"49",x"74",x"4c"),
   834 => (x"ed",x"fd",x"49",x"73"),
   835 => (x"87",x"d6",x"ec",x"87"),
   836 => (x"5c",x"5b",x"5e",x"0e"),
   837 => (x"86",x"f4",x"0e",x"5d"),
   838 => (x"7e",x"c0",x"4a",x"71"),
   839 => (x"d8",x"02",x"9a",x"72"),
   840 => (x"ce",x"f0",x"c3",x"87"),
   841 => (x"c3",x"78",x"c0",x"48"),
   842 => (x"c3",x"48",x"c6",x"f0"),
   843 => (x"78",x"bf",x"ff",x"fc"),
   844 => (x"48",x"ca",x"f0",x"c3"),
   845 => (x"bf",x"fb",x"fc",x"c3"),
   846 => (x"ef",x"f8",x"c3",x"78"),
   847 => (x"c3",x"50",x"c0",x"48"),
   848 => (x"49",x"bf",x"de",x"f8"),
   849 => (x"bf",x"ce",x"f0",x"c3"),
   850 => (x"03",x"aa",x"71",x"4a"),
   851 => (x"72",x"87",x"c0",x"c4"),
   852 => (x"05",x"99",x"cf",x"49"),
   853 => (x"c3",x"87",x"e1",x"c0"),
   854 => (x"c3",x"1e",x"d2",x"f0"),
   855 => (x"49",x"bf",x"c6",x"f0"),
   856 => (x"48",x"c6",x"f0",x"c3"),
   857 => (x"71",x"78",x"a1",x"c1"),
   858 => (x"87",x"fa",x"dc",x"ff"),
   859 => (x"fb",x"c0",x"86",x"c4"),
   860 => (x"f0",x"c3",x"48",x"e4"),
   861 => (x"87",x"cc",x"78",x"d2"),
   862 => (x"bf",x"e4",x"fb",x"c0"),
   863 => (x"80",x"e0",x"c0",x"48"),
   864 => (x"58",x"e8",x"fb",x"c0"),
   865 => (x"bf",x"ce",x"f0",x"c3"),
   866 => (x"c3",x"80",x"c1",x"48"),
   867 => (x"27",x"58",x"d2",x"f0"),
   868 => (x"00",x"00",x"0e",x"e4"),
   869 => (x"4d",x"bf",x"97",x"bf"),
   870 => (x"e2",x"c2",x"02",x"9d"),
   871 => (x"ad",x"e5",x"c3",x"87"),
   872 => (x"87",x"db",x"c2",x"02"),
   873 => (x"bf",x"e4",x"fb",x"c0"),
   874 => (x"49",x"a3",x"cb",x"4b"),
   875 => (x"ac",x"cf",x"4c",x"11"),
   876 => (x"87",x"d2",x"c1",x"05"),
   877 => (x"99",x"df",x"49",x"75"),
   878 => (x"91",x"cd",x"89",x"c1"),
   879 => (x"81",x"e2",x"f8",x"c3"),
   880 => (x"12",x"4a",x"a3",x"c1"),
   881 => (x"4a",x"a3",x"c3",x"51"),
   882 => (x"a3",x"c5",x"51",x"12"),
   883 => (x"c7",x"51",x"12",x"4a"),
   884 => (x"51",x"12",x"4a",x"a3"),
   885 => (x"12",x"4a",x"a3",x"c9"),
   886 => (x"4a",x"a3",x"ce",x"51"),
   887 => (x"a3",x"d0",x"51",x"12"),
   888 => (x"d2",x"51",x"12",x"4a"),
   889 => (x"51",x"12",x"4a",x"a3"),
   890 => (x"12",x"4a",x"a3",x"d4"),
   891 => (x"4a",x"a3",x"d6",x"51"),
   892 => (x"a3",x"d8",x"51",x"12"),
   893 => (x"dc",x"51",x"12",x"4a"),
   894 => (x"51",x"12",x"4a",x"a3"),
   895 => (x"12",x"4a",x"a3",x"de"),
   896 => (x"c0",x"7e",x"c1",x"51"),
   897 => (x"49",x"74",x"87",x"f9"),
   898 => (x"c0",x"05",x"99",x"c8"),
   899 => (x"49",x"74",x"87",x"ea"),
   900 => (x"d0",x"05",x"99",x"d0"),
   901 => (x"02",x"66",x"dc",x"87"),
   902 => (x"73",x"87",x"ca",x"c0"),
   903 => (x"0f",x"66",x"dc",x"49"),
   904 => (x"d3",x"02",x"98",x"70"),
   905 => (x"c0",x"05",x"6e",x"87"),
   906 => (x"f8",x"c3",x"87",x"c6"),
   907 => (x"50",x"c0",x"48",x"e2"),
   908 => (x"bf",x"e4",x"fb",x"c0"),
   909 => (x"87",x"e7",x"c2",x"48"),
   910 => (x"48",x"ef",x"f8",x"c3"),
   911 => (x"c3",x"7e",x"50",x"c0"),
   912 => (x"49",x"bf",x"de",x"f8"),
   913 => (x"bf",x"ce",x"f0",x"c3"),
   914 => (x"04",x"aa",x"71",x"4a"),
   915 => (x"c3",x"87",x"c0",x"fc"),
   916 => (x"05",x"bf",x"ff",x"fc"),
   917 => (x"c3",x"87",x"c8",x"c0"),
   918 => (x"02",x"bf",x"da",x"f8"),
   919 => (x"c0",x"87",x"fe",x"c1"),
   920 => (x"ff",x"48",x"e8",x"fb"),
   921 => (x"ca",x"f0",x"c3",x"78"),
   922 => (x"ff",x"e6",x"49",x"bf"),
   923 => (x"c3",x"49",x"70",x"87"),
   924 => (x"c4",x"59",x"ce",x"f0"),
   925 => (x"f0",x"c3",x"48",x"a6"),
   926 => (x"c3",x"78",x"bf",x"ca"),
   927 => (x"02",x"bf",x"da",x"f8"),
   928 => (x"c4",x"87",x"d8",x"c0"),
   929 => (x"ff",x"cf",x"49",x"66"),
   930 => (x"99",x"f8",x"ff",x"ff"),
   931 => (x"c5",x"c0",x"02",x"a9"),
   932 => (x"c0",x"4d",x"c0",x"87"),
   933 => (x"4d",x"c1",x"87",x"e1"),
   934 => (x"c4",x"87",x"dc",x"c0"),
   935 => (x"ff",x"cf",x"49",x"66"),
   936 => (x"02",x"a9",x"99",x"f8"),
   937 => (x"c8",x"87",x"c8",x"c0"),
   938 => (x"78",x"c0",x"48",x"a6"),
   939 => (x"c8",x"87",x"c5",x"c0"),
   940 => (x"78",x"c1",x"48",x"a6"),
   941 => (x"75",x"4d",x"66",x"c8"),
   942 => (x"e0",x"c0",x"05",x"9d"),
   943 => (x"49",x"66",x"c4",x"87"),
   944 => (x"f8",x"c3",x"89",x"c2"),
   945 => (x"91",x"4a",x"bf",x"d2"),
   946 => (x"bf",x"eb",x"fc",x"c3"),
   947 => (x"c6",x"f0",x"c3",x"4a"),
   948 => (x"78",x"a1",x"72",x"48"),
   949 => (x"48",x"ce",x"f0",x"c3"),
   950 => (x"e2",x"f9",x"78",x"c0"),
   951 => (x"f4",x"48",x"c0",x"87"),
   952 => (x"87",x"c0",x"e5",x"8e"),
   953 => (x"00",x"00",x"00",x"00"),
   954 => (x"ff",x"ff",x"ff",x"ff"),
   955 => (x"00",x"00",x"0e",x"f4"),
   956 => (x"00",x"00",x"0e",x"fd"),
   957 => (x"33",x"54",x"41",x"46"),
   958 => (x"20",x"20",x"20",x"32"),
   959 => (x"54",x"41",x"46",x"00"),
   960 => (x"20",x"20",x"36",x"31"),
   961 => (x"ff",x"1e",x"00",x"20"),
   962 => (x"ff",x"c3",x"48",x"d4"),
   963 => (x"26",x"48",x"68",x"78"),
   964 => (x"d4",x"ff",x"1e",x"4f"),
   965 => (x"78",x"ff",x"c3",x"48"),
   966 => (x"c8",x"48",x"d0",x"ff"),
   967 => (x"d4",x"ff",x"78",x"e1"),
   968 => (x"c3",x"78",x"d4",x"48"),
   969 => (x"ff",x"48",x"c3",x"fd"),
   970 => (x"26",x"50",x"bf",x"d4"),
   971 => (x"d0",x"ff",x"1e",x"4f"),
   972 => (x"78",x"e0",x"c0",x"48"),
   973 => (x"ff",x"1e",x"4f",x"26"),
   974 => (x"49",x"70",x"87",x"cc"),
   975 => (x"87",x"c6",x"02",x"99"),
   976 => (x"05",x"a9",x"fb",x"c0"),
   977 => (x"48",x"71",x"87",x"f1"),
   978 => (x"5e",x"0e",x"4f",x"26"),
   979 => (x"71",x"0e",x"5c",x"5b"),
   980 => (x"fe",x"4c",x"c0",x"4b"),
   981 => (x"49",x"70",x"87",x"f0"),
   982 => (x"f9",x"c0",x"02",x"99"),
   983 => (x"a9",x"ec",x"c0",x"87"),
   984 => (x"87",x"f2",x"c0",x"02"),
   985 => (x"02",x"a9",x"fb",x"c0"),
   986 => (x"cc",x"87",x"eb",x"c0"),
   987 => (x"03",x"ac",x"b7",x"66"),
   988 => (x"66",x"d0",x"87",x"c7"),
   989 => (x"71",x"87",x"c2",x"02"),
   990 => (x"02",x"99",x"71",x"53"),
   991 => (x"84",x"c1",x"87",x"c2"),
   992 => (x"70",x"87",x"c3",x"fe"),
   993 => (x"cd",x"02",x"99",x"49"),
   994 => (x"a9",x"ec",x"c0",x"87"),
   995 => (x"c0",x"87",x"c7",x"02"),
   996 => (x"ff",x"05",x"a9",x"fb"),
   997 => (x"66",x"d0",x"87",x"d5"),
   998 => (x"c0",x"87",x"c3",x"02"),
   999 => (x"ec",x"c0",x"7b",x"97"),
  1000 => (x"87",x"c4",x"05",x"a9"),
  1001 => (x"87",x"c5",x"4a",x"74"),
  1002 => (x"0a",x"c0",x"4a",x"74"),
  1003 => (x"c2",x"48",x"72",x"8a"),
  1004 => (x"26",x"4d",x"26",x"87"),
  1005 => (x"26",x"4b",x"26",x"4c"),
  1006 => (x"c9",x"fd",x"1e",x"4f"),
  1007 => (x"c0",x"49",x"70",x"87"),
  1008 => (x"04",x"a9",x"b7",x"f0"),
  1009 => (x"f9",x"c0",x"87",x"ca"),
  1010 => (x"c3",x"01",x"a9",x"b7"),
  1011 => (x"89",x"f0",x"c0",x"87"),
  1012 => (x"a9",x"b7",x"c1",x"c1"),
  1013 => (x"c1",x"87",x"ca",x"04"),
  1014 => (x"01",x"a9",x"b7",x"da"),
  1015 => (x"f7",x"c0",x"87",x"c3"),
  1016 => (x"26",x"48",x"71",x"89"),
  1017 => (x"5b",x"5e",x"0e",x"4f"),
  1018 => (x"4c",x"71",x"0e",x"5c"),
  1019 => (x"c1",x"87",x"e2",x"fc"),
  1020 => (x"1e",x"66",x"d0",x"1e"),
  1021 => (x"d1",x"fd",x"49",x"74"),
  1022 => (x"70",x"86",x"c8",x"87"),
  1023 => (x"87",x"ed",x"fc",x"4b"),
  1024 => (x"03",x"ab",x"b7",x"c0"),
  1025 => (x"8b",x"0b",x"87",x"c2"),
  1026 => (x"ab",x"b7",x"66",x"cc"),
  1027 => (x"74",x"87",x"cf",x"03"),
  1028 => (x"83",x"c1",x"49",x"a3"),
  1029 => (x"cc",x"51",x"e0",x"c0"),
  1030 => (x"04",x"ab",x"b7",x"66"),
  1031 => (x"a3",x"74",x"87",x"f1"),
  1032 => (x"fe",x"51",x"c0",x"49"),
  1033 => (x"5e",x"0e",x"87",x"cd"),
  1034 => (x"71",x"0e",x"5c",x"5b"),
  1035 => (x"4c",x"d4",x"ff",x"4a"),
  1036 => (x"ea",x"c0",x"49",x"72"),
  1037 => (x"9b",x"4b",x"70",x"87"),
  1038 => (x"c1",x"87",x"c2",x"02"),
  1039 => (x"48",x"d0",x"ff",x"8b"),
  1040 => (x"c1",x"78",x"c5",x"c8"),
  1041 => (x"49",x"73",x"7c",x"d5"),
  1042 => (x"cf",x"c3",x"31",x"c6"),
  1043 => (x"4a",x"bf",x"97",x"da"),
  1044 => (x"70",x"b0",x"71",x"48"),
  1045 => (x"48",x"d0",x"ff",x"7c"),
  1046 => (x"48",x"73",x"78",x"c4"),
  1047 => (x"0e",x"87",x"d4",x"fd"),
  1048 => (x"5d",x"5c",x"5b",x"5e"),
  1049 => (x"71",x"86",x"f8",x"0e"),
  1050 => (x"fa",x"7e",x"c0",x"4c"),
  1051 => (x"4b",x"c0",x"87",x"e3"),
  1052 => (x"97",x"cc",x"c4",x"c1"),
  1053 => (x"a9",x"c0",x"49",x"bf"),
  1054 => (x"fa",x"87",x"cf",x"04"),
  1055 => (x"83",x"c1",x"87",x"f8"),
  1056 => (x"97",x"cc",x"c4",x"c1"),
  1057 => (x"06",x"ab",x"49",x"bf"),
  1058 => (x"c4",x"c1",x"87",x"f1"),
  1059 => (x"02",x"bf",x"97",x"cc"),
  1060 => (x"f1",x"f9",x"87",x"cf"),
  1061 => (x"99",x"49",x"70",x"87"),
  1062 => (x"c0",x"87",x"c6",x"02"),
  1063 => (x"f1",x"05",x"a9",x"ec"),
  1064 => (x"f9",x"4b",x"c0",x"87"),
  1065 => (x"4d",x"70",x"87",x"e0"),
  1066 => (x"c8",x"87",x"db",x"f9"),
  1067 => (x"d5",x"f9",x"58",x"a6"),
  1068 => (x"c1",x"4a",x"70",x"87"),
  1069 => (x"49",x"a4",x"c8",x"83"),
  1070 => (x"ad",x"49",x"69",x"97"),
  1071 => (x"c0",x"87",x"c7",x"02"),
  1072 => (x"c0",x"05",x"ad",x"ff"),
  1073 => (x"a4",x"c9",x"87",x"e7"),
  1074 => (x"49",x"69",x"97",x"49"),
  1075 => (x"02",x"a9",x"66",x"c4"),
  1076 => (x"c0",x"48",x"87",x"c7"),
  1077 => (x"d4",x"05",x"a8",x"ff"),
  1078 => (x"49",x"a4",x"ca",x"87"),
  1079 => (x"aa",x"49",x"69",x"97"),
  1080 => (x"c0",x"87",x"c6",x"02"),
  1081 => (x"c4",x"05",x"aa",x"ff"),
  1082 => (x"d0",x"7e",x"c1",x"87"),
  1083 => (x"ad",x"ec",x"c0",x"87"),
  1084 => (x"c0",x"87",x"c6",x"02"),
  1085 => (x"c4",x"05",x"ad",x"fb"),
  1086 => (x"c1",x"4b",x"c0",x"87"),
  1087 => (x"fe",x"02",x"6e",x"7e"),
  1088 => (x"e8",x"f8",x"87",x"e1"),
  1089 => (x"f8",x"48",x"73",x"87"),
  1090 => (x"87",x"e5",x"fa",x"8e"),
  1091 => (x"5b",x"5e",x"0e",x"00"),
  1092 => (x"1e",x"0e",x"5d",x"5c"),
  1093 => (x"4c",x"c0",x"4b",x"71"),
  1094 => (x"c0",x"04",x"ab",x"4d"),
  1095 => (x"c1",x"c1",x"87",x"e8"),
  1096 => (x"9d",x"75",x"1e",x"df"),
  1097 => (x"c0",x"87",x"c4",x"02"),
  1098 => (x"c1",x"87",x"c2",x"4a"),
  1099 => (x"ef",x"49",x"72",x"4a"),
  1100 => (x"86",x"c4",x"87",x"de"),
  1101 => (x"84",x"c1",x"7e",x"70"),
  1102 => (x"87",x"c2",x"05",x"6e"),
  1103 => (x"85",x"c1",x"4c",x"73"),
  1104 => (x"ff",x"06",x"ac",x"73"),
  1105 => (x"48",x"6e",x"87",x"d8"),
  1106 => (x"26",x"4d",x"26",x"26"),
  1107 => (x"26",x"4b",x"26",x"4c"),
  1108 => (x"5b",x"5e",x"0e",x"4f"),
  1109 => (x"1e",x"0e",x"5d",x"5c"),
  1110 => (x"de",x"49",x"4c",x"71"),
  1111 => (x"dd",x"fd",x"c3",x"91"),
  1112 => (x"97",x"85",x"71",x"4d"),
  1113 => (x"dd",x"c1",x"02",x"6d"),
  1114 => (x"c8",x"fd",x"c3",x"87"),
  1115 => (x"82",x"74",x"4a",x"bf"),
  1116 => (x"d8",x"fe",x"49",x"72"),
  1117 => (x"6e",x"7e",x"70",x"87"),
  1118 => (x"87",x"f3",x"c0",x"02"),
  1119 => (x"4b",x"d0",x"fd",x"c3"),
  1120 => (x"49",x"cb",x"4a",x"6e"),
  1121 => (x"87",x"de",x"fd",x"fe"),
  1122 => (x"93",x"cb",x"4b",x"74"),
  1123 => (x"83",x"d7",x"e9",x"c1"),
  1124 => (x"c7",x"c1",x"83",x"c4"),
  1125 => (x"49",x"74",x"7b",x"ca"),
  1126 => (x"87",x"e5",x"c4",x"c1"),
  1127 => (x"fd",x"c3",x"7b",x"75"),
  1128 => (x"49",x"bf",x"97",x"dc"),
  1129 => (x"d0",x"fd",x"c3",x"1e"),
  1130 => (x"c0",x"da",x"c2",x"49"),
  1131 => (x"74",x"86",x"c4",x"87"),
  1132 => (x"cc",x"c4",x"c1",x"49"),
  1133 => (x"c1",x"49",x"c0",x"87"),
  1134 => (x"c3",x"87",x"eb",x"c5"),
  1135 => (x"c0",x"48",x"c4",x"fd"),
  1136 => (x"dd",x"49",x"c1",x"78"),
  1137 => (x"fd",x"26",x"87",x"d1"),
  1138 => (x"6f",x"4c",x"87",x"ff"),
  1139 => (x"6e",x"69",x"64",x"61"),
  1140 => (x"2e",x"2e",x"2e",x"67"),
  1141 => (x"5b",x"5e",x"0e",x"00"),
  1142 => (x"4b",x"71",x"0e",x"5c"),
  1143 => (x"c8",x"fd",x"c3",x"4a"),
  1144 => (x"49",x"72",x"82",x"bf"),
  1145 => (x"70",x"87",x"e6",x"fc"),
  1146 => (x"c4",x"02",x"9c",x"4c"),
  1147 => (x"e7",x"eb",x"49",x"87"),
  1148 => (x"c8",x"fd",x"c3",x"87"),
  1149 => (x"c1",x"78",x"c0",x"48"),
  1150 => (x"87",x"db",x"dc",x"49"),
  1151 => (x"0e",x"87",x"cc",x"fd"),
  1152 => (x"5d",x"5c",x"5b",x"5e"),
  1153 => (x"c3",x"86",x"f4",x"0e"),
  1154 => (x"c0",x"4d",x"d2",x"f0"),
  1155 => (x"48",x"a6",x"c4",x"4c"),
  1156 => (x"fd",x"c3",x"78",x"c0"),
  1157 => (x"c0",x"49",x"bf",x"c8"),
  1158 => (x"c1",x"c1",x"06",x"a9"),
  1159 => (x"d2",x"f0",x"c3",x"87"),
  1160 => (x"c0",x"02",x"98",x"48"),
  1161 => (x"c1",x"c1",x"87",x"f8"),
  1162 => (x"66",x"c8",x"1e",x"df"),
  1163 => (x"c4",x"87",x"c7",x"02"),
  1164 => (x"78",x"c0",x"48",x"a6"),
  1165 => (x"a6",x"c4",x"87",x"c5"),
  1166 => (x"c4",x"78",x"c1",x"48"),
  1167 => (x"cf",x"eb",x"49",x"66"),
  1168 => (x"70",x"86",x"c4",x"87"),
  1169 => (x"c4",x"84",x"c1",x"4d"),
  1170 => (x"80",x"c1",x"48",x"66"),
  1171 => (x"c3",x"58",x"a6",x"c8"),
  1172 => (x"49",x"bf",x"c8",x"fd"),
  1173 => (x"87",x"c6",x"03",x"ac"),
  1174 => (x"ff",x"05",x"9d",x"75"),
  1175 => (x"4c",x"c0",x"87",x"c8"),
  1176 => (x"c3",x"02",x"9d",x"75"),
  1177 => (x"c1",x"c1",x"87",x"e0"),
  1178 => (x"66",x"c8",x"1e",x"df"),
  1179 => (x"cc",x"87",x"c7",x"02"),
  1180 => (x"78",x"c0",x"48",x"a6"),
  1181 => (x"a6",x"cc",x"87",x"c5"),
  1182 => (x"cc",x"78",x"c1",x"48"),
  1183 => (x"cf",x"ea",x"49",x"66"),
  1184 => (x"70",x"86",x"c4",x"87"),
  1185 => (x"c2",x"02",x"6e",x"7e"),
  1186 => (x"49",x"6e",x"87",x"e9"),
  1187 => (x"69",x"97",x"81",x"cb"),
  1188 => (x"02",x"99",x"d0",x"49"),
  1189 => (x"c1",x"87",x"d6",x"c1"),
  1190 => (x"74",x"4a",x"d5",x"c7"),
  1191 => (x"c1",x"91",x"cb",x"49"),
  1192 => (x"72",x"81",x"d7",x"e9"),
  1193 => (x"c3",x"81",x"c8",x"79"),
  1194 => (x"49",x"74",x"51",x"ff"),
  1195 => (x"fd",x"c3",x"91",x"de"),
  1196 => (x"85",x"71",x"4d",x"dd"),
  1197 => (x"7d",x"97",x"c1",x"c2"),
  1198 => (x"c0",x"49",x"a5",x"c1"),
  1199 => (x"f8",x"c3",x"51",x"e0"),
  1200 => (x"02",x"bf",x"97",x"e2"),
  1201 => (x"84",x"c1",x"87",x"d2"),
  1202 => (x"c3",x"4b",x"a5",x"c2"),
  1203 => (x"db",x"4a",x"e2",x"f8"),
  1204 => (x"d1",x"f8",x"fe",x"49"),
  1205 => (x"87",x"db",x"c1",x"87"),
  1206 => (x"c0",x"49",x"a5",x"cd"),
  1207 => (x"c2",x"84",x"c1",x"51"),
  1208 => (x"4a",x"6e",x"4b",x"a5"),
  1209 => (x"f7",x"fe",x"49",x"cb"),
  1210 => (x"c6",x"c1",x"87",x"fc"),
  1211 => (x"d1",x"c5",x"c1",x"87"),
  1212 => (x"cb",x"49",x"74",x"4a"),
  1213 => (x"d7",x"e9",x"c1",x"91"),
  1214 => (x"c3",x"79",x"72",x"81"),
  1215 => (x"bf",x"97",x"e2",x"f8"),
  1216 => (x"74",x"87",x"d8",x"02"),
  1217 => (x"c1",x"91",x"de",x"49"),
  1218 => (x"dd",x"fd",x"c3",x"84"),
  1219 => (x"c3",x"83",x"71",x"4b"),
  1220 => (x"dd",x"4a",x"e2",x"f8"),
  1221 => (x"cd",x"f7",x"fe",x"49"),
  1222 => (x"74",x"87",x"d8",x"87"),
  1223 => (x"c3",x"93",x"de",x"4b"),
  1224 => (x"cb",x"83",x"dd",x"fd"),
  1225 => (x"51",x"c0",x"49",x"a3"),
  1226 => (x"6e",x"73",x"84",x"c1"),
  1227 => (x"fe",x"49",x"cb",x"4a"),
  1228 => (x"c4",x"87",x"f3",x"f6"),
  1229 => (x"80",x"c1",x"48",x"66"),
  1230 => (x"c7",x"58",x"a6",x"c8"),
  1231 => (x"c5",x"c0",x"03",x"ac"),
  1232 => (x"fc",x"05",x"6e",x"87"),
  1233 => (x"48",x"74",x"87",x"e0"),
  1234 => (x"fc",x"f7",x"8e",x"f4"),
  1235 => (x"1e",x"73",x"1e",x"87"),
  1236 => (x"cb",x"49",x"4b",x"71"),
  1237 => (x"d7",x"e9",x"c1",x"91"),
  1238 => (x"4a",x"a1",x"c8",x"81"),
  1239 => (x"48",x"da",x"cf",x"c3"),
  1240 => (x"a1",x"c9",x"50",x"12"),
  1241 => (x"cc",x"c4",x"c1",x"4a"),
  1242 => (x"ca",x"50",x"12",x"48"),
  1243 => (x"dc",x"fd",x"c3",x"81"),
  1244 => (x"c3",x"50",x"11",x"48"),
  1245 => (x"bf",x"97",x"dc",x"fd"),
  1246 => (x"49",x"c0",x"1e",x"49"),
  1247 => (x"87",x"ed",x"d2",x"c2"),
  1248 => (x"48",x"c4",x"fd",x"c3"),
  1249 => (x"49",x"c1",x"78",x"de"),
  1250 => (x"26",x"87",x"cc",x"d6"),
  1251 => (x"1e",x"87",x"fe",x"f6"),
  1252 => (x"cb",x"49",x"4a",x"71"),
  1253 => (x"d7",x"e9",x"c1",x"91"),
  1254 => (x"11",x"81",x"c8",x"81"),
  1255 => (x"c8",x"fd",x"c3",x"48"),
  1256 => (x"c8",x"fd",x"c3",x"58"),
  1257 => (x"c1",x"78",x"c0",x"48"),
  1258 => (x"87",x"eb",x"d5",x"49"),
  1259 => (x"c0",x"1e",x"4f",x"26"),
  1260 => (x"f1",x"fd",x"c0",x"49"),
  1261 => (x"1e",x"4f",x"26",x"87"),
  1262 => (x"d2",x"02",x"99",x"71"),
  1263 => (x"ec",x"ea",x"c1",x"87"),
  1264 => (x"f7",x"50",x"c0",x"48"),
  1265 => (x"cf",x"ce",x"c1",x"80"),
  1266 => (x"d0",x"e9",x"c1",x"40"),
  1267 => (x"c1",x"87",x"ce",x"78"),
  1268 => (x"c1",x"48",x"e8",x"ea"),
  1269 => (x"fc",x"78",x"c9",x"e9"),
  1270 => (x"ee",x"ce",x"c1",x"80"),
  1271 => (x"0e",x"4f",x"26",x"78"),
  1272 => (x"0e",x"5c",x"5b",x"5e"),
  1273 => (x"cb",x"4a",x"4c",x"71"),
  1274 => (x"d7",x"e9",x"c1",x"92"),
  1275 => (x"49",x"a2",x"c8",x"82"),
  1276 => (x"97",x"4b",x"a2",x"c9"),
  1277 => (x"97",x"1e",x"4b",x"6b"),
  1278 => (x"ca",x"1e",x"49",x"69"),
  1279 => (x"c0",x"49",x"12",x"82"),
  1280 => (x"c0",x"87",x"ec",x"e8"),
  1281 => (x"87",x"cf",x"d4",x"49"),
  1282 => (x"fa",x"c0",x"49",x"74"),
  1283 => (x"8e",x"f8",x"87",x"f3"),
  1284 => (x"1e",x"87",x"f8",x"f4"),
  1285 => (x"4b",x"71",x"1e",x"73"),
  1286 => (x"87",x"c3",x"ff",x"49"),
  1287 => (x"fe",x"fe",x"49",x"73"),
  1288 => (x"c0",x"49",x"c0",x"87"),
  1289 => (x"f4",x"87",x"ff",x"fb"),
  1290 => (x"73",x"1e",x"87",x"e3"),
  1291 => (x"c6",x"4b",x"71",x"1e"),
  1292 => (x"db",x"02",x"4a",x"a3"),
  1293 => (x"02",x"8a",x"c1",x"87"),
  1294 => (x"02",x"8a",x"87",x"d6"),
  1295 => (x"8a",x"87",x"da",x"c1"),
  1296 => (x"87",x"fc",x"c0",x"02"),
  1297 => (x"e1",x"c0",x"02",x"8a"),
  1298 => (x"cb",x"02",x"8a",x"87"),
  1299 => (x"87",x"db",x"c1",x"87"),
  1300 => (x"fa",x"fc",x"49",x"c7"),
  1301 => (x"87",x"de",x"c1",x"87"),
  1302 => (x"bf",x"c8",x"fd",x"c3"),
  1303 => (x"87",x"cb",x"c1",x"02"),
  1304 => (x"c3",x"88",x"c1",x"48"),
  1305 => (x"c1",x"58",x"cc",x"fd"),
  1306 => (x"fd",x"c3",x"87",x"c1"),
  1307 => (x"c0",x"02",x"bf",x"cc"),
  1308 => (x"fd",x"c3",x"87",x"f9"),
  1309 => (x"c1",x"48",x"bf",x"c8"),
  1310 => (x"cc",x"fd",x"c3",x"80"),
  1311 => (x"87",x"eb",x"c0",x"58"),
  1312 => (x"bf",x"c8",x"fd",x"c3"),
  1313 => (x"c3",x"89",x"c6",x"49"),
  1314 => (x"c0",x"59",x"cc",x"fd"),
  1315 => (x"da",x"03",x"a9",x"b7"),
  1316 => (x"c8",x"fd",x"c3",x"87"),
  1317 => (x"d2",x"78",x"c0",x"48"),
  1318 => (x"cc",x"fd",x"c3",x"87"),
  1319 => (x"87",x"cb",x"02",x"bf"),
  1320 => (x"bf",x"c8",x"fd",x"c3"),
  1321 => (x"c3",x"80",x"c6",x"48"),
  1322 => (x"c0",x"58",x"cc",x"fd"),
  1323 => (x"87",x"e7",x"d1",x"49"),
  1324 => (x"f8",x"c0",x"49",x"73"),
  1325 => (x"d4",x"f2",x"87",x"cb"),
  1326 => (x"5b",x"5e",x"0e",x"87"),
  1327 => (x"4c",x"71",x"0e",x"5c"),
  1328 => (x"74",x"1e",x"66",x"cc"),
  1329 => (x"c1",x"93",x"cb",x"4b"),
  1330 => (x"c4",x"83",x"d7",x"e9"),
  1331 => (x"49",x"6a",x"4a",x"a3"),
  1332 => (x"87",x"e2",x"f0",x"fe"),
  1333 => (x"7b",x"cd",x"cd",x"c1"),
  1334 => (x"d4",x"49",x"a3",x"c8"),
  1335 => (x"a3",x"c9",x"51",x"66"),
  1336 => (x"51",x"66",x"d8",x"49"),
  1337 => (x"dc",x"49",x"a3",x"ca"),
  1338 => (x"f1",x"26",x"51",x"66"),
  1339 => (x"5e",x"0e",x"87",x"dd"),
  1340 => (x"0e",x"5d",x"5c",x"5b"),
  1341 => (x"d8",x"86",x"d0",x"ff"),
  1342 => (x"a6",x"c4",x"59",x"a6"),
  1343 => (x"c4",x"78",x"c0",x"48"),
  1344 => (x"66",x"c4",x"c1",x"80"),
  1345 => (x"c1",x"80",x"c4",x"78"),
  1346 => (x"c1",x"80",x"c4",x"78"),
  1347 => (x"cc",x"fd",x"c3",x"78"),
  1348 => (x"c3",x"78",x"c1",x"48"),
  1349 => (x"48",x"bf",x"c4",x"fd"),
  1350 => (x"cb",x"05",x"a8",x"de"),
  1351 => (x"87",x"df",x"f3",x"87"),
  1352 => (x"a6",x"c8",x"49",x"70"),
  1353 => (x"87",x"f8",x"ce",x"59"),
  1354 => (x"e8",x"87",x"e6",x"e7"),
  1355 => (x"d5",x"e7",x"87",x"c8"),
  1356 => (x"c0",x"4c",x"70",x"87"),
  1357 => (x"c1",x"02",x"ac",x"fb"),
  1358 => (x"66",x"d4",x"87",x"d0"),
  1359 => (x"87",x"c2",x"c1",x"05"),
  1360 => (x"c1",x"1e",x"1e",x"c0"),
  1361 => (x"fa",x"ea",x"c1",x"1e"),
  1362 => (x"fd",x"49",x"c0",x"1e"),
  1363 => (x"d0",x"c1",x"87",x"eb"),
  1364 => (x"82",x"c4",x"4a",x"66"),
  1365 => (x"81",x"c7",x"49",x"6a"),
  1366 => (x"1e",x"c1",x"51",x"74"),
  1367 => (x"49",x"6a",x"1e",x"d8"),
  1368 => (x"e5",x"e7",x"81",x"c8"),
  1369 => (x"c1",x"86",x"d8",x"87"),
  1370 => (x"c0",x"48",x"66",x"c4"),
  1371 => (x"87",x"c7",x"01",x"a8"),
  1372 => (x"c1",x"48",x"a6",x"c4"),
  1373 => (x"c1",x"87",x"ce",x"78"),
  1374 => (x"c1",x"48",x"66",x"c4"),
  1375 => (x"58",x"a6",x"cc",x"88"),
  1376 => (x"f1",x"e6",x"87",x"c3"),
  1377 => (x"48",x"a6",x"cc",x"87"),
  1378 => (x"9c",x"74",x"78",x"c2"),
  1379 => (x"87",x"cc",x"cd",x"02"),
  1380 => (x"c1",x"48",x"66",x"c4"),
  1381 => (x"03",x"a8",x"66",x"c8"),
  1382 => (x"d8",x"87",x"c1",x"cd"),
  1383 => (x"78",x"c0",x"48",x"a6"),
  1384 => (x"70",x"87",x"e3",x"e5"),
  1385 => (x"ac",x"d0",x"c1",x"4c"),
  1386 => (x"87",x"d6",x"c2",x"05"),
  1387 => (x"e8",x"7e",x"66",x"d8"),
  1388 => (x"49",x"70",x"87",x"c7"),
  1389 => (x"e5",x"59",x"a6",x"dc"),
  1390 => (x"4c",x"70",x"87",x"cc"),
  1391 => (x"05",x"ac",x"ec",x"c0"),
  1392 => (x"c4",x"87",x"ea",x"c1"),
  1393 => (x"91",x"cb",x"49",x"66"),
  1394 => (x"81",x"66",x"c0",x"c1"),
  1395 => (x"6a",x"4a",x"a1",x"c4"),
  1396 => (x"4a",x"a1",x"c8",x"4d"),
  1397 => (x"c1",x"52",x"66",x"d8"),
  1398 => (x"e4",x"79",x"cf",x"ce"),
  1399 => (x"4c",x"70",x"87",x"e8"),
  1400 => (x"87",x"d8",x"02",x"9c"),
  1401 => (x"02",x"ac",x"fb",x"c0"),
  1402 => (x"55",x"74",x"87",x"d2"),
  1403 => (x"70",x"87",x"d7",x"e4"),
  1404 => (x"c7",x"02",x"9c",x"4c"),
  1405 => (x"ac",x"fb",x"c0",x"87"),
  1406 => (x"87",x"ee",x"ff",x"05"),
  1407 => (x"c2",x"55",x"e0",x"c0"),
  1408 => (x"97",x"c0",x"55",x"c1"),
  1409 => (x"49",x"66",x"d4",x"7d"),
  1410 => (x"db",x"05",x"a9",x"6e"),
  1411 => (x"48",x"66",x"c4",x"87"),
  1412 => (x"04",x"a8",x"66",x"c8"),
  1413 => (x"66",x"c4",x"87",x"ca"),
  1414 => (x"c8",x"80",x"c1",x"48"),
  1415 => (x"87",x"c8",x"58",x"a6"),
  1416 => (x"c1",x"48",x"66",x"c8"),
  1417 => (x"58",x"a6",x"cc",x"88"),
  1418 => (x"70",x"87",x"db",x"e3"),
  1419 => (x"ac",x"d0",x"c1",x"4c"),
  1420 => (x"d0",x"87",x"c8",x"05"),
  1421 => (x"80",x"c1",x"48",x"66"),
  1422 => (x"c1",x"58",x"a6",x"d4"),
  1423 => (x"fd",x"02",x"ac",x"d0"),
  1424 => (x"a6",x"dc",x"87",x"ea"),
  1425 => (x"78",x"66",x"d4",x"48"),
  1426 => (x"dc",x"48",x"66",x"d8"),
  1427 => (x"c9",x"05",x"a8",x"66"),
  1428 => (x"e0",x"c0",x"87",x"dc"),
  1429 => (x"f0",x"c0",x"48",x"a6"),
  1430 => (x"cc",x"80",x"c4",x"78"),
  1431 => (x"80",x"c4",x"78",x"66"),
  1432 => (x"74",x"7e",x"78",x"c0"),
  1433 => (x"88",x"fb",x"c0",x"48"),
  1434 => (x"58",x"a6",x"f0",x"c0"),
  1435 => (x"c8",x"02",x"98",x"70"),
  1436 => (x"cb",x"48",x"87",x"d7"),
  1437 => (x"a6",x"f0",x"c0",x"88"),
  1438 => (x"02",x"98",x"70",x"58"),
  1439 => (x"48",x"87",x"e9",x"c0"),
  1440 => (x"f0",x"c0",x"88",x"c9"),
  1441 => (x"98",x"70",x"58",x"a6"),
  1442 => (x"87",x"e1",x"c3",x"02"),
  1443 => (x"c0",x"88",x"c4",x"48"),
  1444 => (x"70",x"58",x"a6",x"f0"),
  1445 => (x"87",x"d6",x"02",x"98"),
  1446 => (x"c0",x"88",x"c1",x"48"),
  1447 => (x"70",x"58",x"a6",x"f0"),
  1448 => (x"c8",x"c3",x"02",x"98"),
  1449 => (x"87",x"db",x"c7",x"87"),
  1450 => (x"48",x"a6",x"e0",x"c0"),
  1451 => (x"66",x"cc",x"78",x"c0"),
  1452 => (x"d0",x"80",x"c1",x"48"),
  1453 => (x"cd",x"e1",x"58",x"a6"),
  1454 => (x"c0",x"4c",x"70",x"87"),
  1455 => (x"d5",x"02",x"ac",x"ec"),
  1456 => (x"66",x"e0",x"c0",x"87"),
  1457 => (x"c0",x"87",x"c6",x"02"),
  1458 => (x"c9",x"5c",x"a6",x"e4"),
  1459 => (x"c0",x"48",x"74",x"87"),
  1460 => (x"e8",x"c0",x"88",x"f0"),
  1461 => (x"ec",x"c0",x"58",x"a6"),
  1462 => (x"87",x"cc",x"02",x"ac"),
  1463 => (x"70",x"87",x"e7",x"e0"),
  1464 => (x"ac",x"ec",x"c0",x"4c"),
  1465 => (x"87",x"f4",x"ff",x"05"),
  1466 => (x"1e",x"66",x"e0",x"c0"),
  1467 => (x"1e",x"49",x"66",x"d4"),
  1468 => (x"1e",x"66",x"ec",x"c0"),
  1469 => (x"1e",x"fa",x"ea",x"c1"),
  1470 => (x"f6",x"49",x"66",x"d4"),
  1471 => (x"1e",x"c0",x"87",x"fb"),
  1472 => (x"66",x"dc",x"1e",x"ca"),
  1473 => (x"c1",x"91",x"cb",x"49"),
  1474 => (x"d8",x"81",x"66",x"d8"),
  1475 => (x"a1",x"c4",x"48",x"a6"),
  1476 => (x"bf",x"66",x"d8",x"78"),
  1477 => (x"87",x"f2",x"e0",x"49"),
  1478 => (x"b7",x"c0",x"86",x"d8"),
  1479 => (x"c7",x"c1",x"06",x"a8"),
  1480 => (x"de",x"1e",x"c1",x"87"),
  1481 => (x"bf",x"66",x"c8",x"1e"),
  1482 => (x"87",x"de",x"e0",x"49"),
  1483 => (x"49",x"70",x"86",x"c8"),
  1484 => (x"88",x"08",x"c0",x"48"),
  1485 => (x"58",x"a6",x"e4",x"c0"),
  1486 => (x"06",x"a8",x"b7",x"c0"),
  1487 => (x"c0",x"87",x"e9",x"c0"),
  1488 => (x"dd",x"48",x"66",x"e0"),
  1489 => (x"df",x"03",x"a8",x"b7"),
  1490 => (x"49",x"bf",x"6e",x"87"),
  1491 => (x"81",x"66",x"e0",x"c0"),
  1492 => (x"66",x"51",x"e0",x"c0"),
  1493 => (x"6e",x"81",x"c1",x"49"),
  1494 => (x"c1",x"c2",x"81",x"bf"),
  1495 => (x"66",x"e0",x"c0",x"51"),
  1496 => (x"6e",x"81",x"c2",x"49"),
  1497 => (x"51",x"c0",x"81",x"bf"),
  1498 => (x"dc",x"c4",x"7e",x"c1"),
  1499 => (x"87",x"c9",x"e1",x"87"),
  1500 => (x"58",x"a6",x"e4",x"c0"),
  1501 => (x"c0",x"87",x"c2",x"e1"),
  1502 => (x"c0",x"58",x"a6",x"e8"),
  1503 => (x"c0",x"05",x"a8",x"ec"),
  1504 => (x"e4",x"c0",x"87",x"cb"),
  1505 => (x"e0",x"c0",x"48",x"a6"),
  1506 => (x"c4",x"c0",x"78",x"66"),
  1507 => (x"f5",x"dd",x"ff",x"87"),
  1508 => (x"49",x"66",x"c4",x"87"),
  1509 => (x"c0",x"c1",x"91",x"cb"),
  1510 => (x"80",x"71",x"48",x"66"),
  1511 => (x"4a",x"6e",x"7e",x"70"),
  1512 => (x"49",x"6e",x"82",x"c8"),
  1513 => (x"e0",x"c0",x"81",x"ca"),
  1514 => (x"e4",x"c0",x"51",x"66"),
  1515 => (x"81",x"c1",x"49",x"66"),
  1516 => (x"89",x"66",x"e0",x"c0"),
  1517 => (x"30",x"71",x"48",x"c1"),
  1518 => (x"89",x"c1",x"49",x"70"),
  1519 => (x"c4",x"7a",x"97",x"71"),
  1520 => (x"49",x"bf",x"f9",x"c0"),
  1521 => (x"29",x"66",x"e0",x"c0"),
  1522 => (x"48",x"4a",x"6a",x"97"),
  1523 => (x"f0",x"c0",x"98",x"71"),
  1524 => (x"49",x"6e",x"58",x"a6"),
  1525 => (x"4d",x"69",x"81",x"c4"),
  1526 => (x"d8",x"48",x"66",x"dc"),
  1527 => (x"c0",x"02",x"a8",x"66"),
  1528 => (x"a6",x"d8",x"87",x"c8"),
  1529 => (x"c0",x"78",x"c0",x"48"),
  1530 => (x"a6",x"d8",x"87",x"c5"),
  1531 => (x"d8",x"78",x"c1",x"48"),
  1532 => (x"e0",x"c0",x"1e",x"66"),
  1533 => (x"ff",x"49",x"75",x"1e"),
  1534 => (x"c8",x"87",x"cf",x"dd"),
  1535 => (x"c0",x"4c",x"70",x"86"),
  1536 => (x"c1",x"06",x"ac",x"b7"),
  1537 => (x"85",x"74",x"87",x"d4"),
  1538 => (x"74",x"49",x"e0",x"c0"),
  1539 => (x"c1",x"4b",x"75",x"89"),
  1540 => (x"71",x"4a",x"d4",x"e4"),
  1541 => (x"87",x"ce",x"e3",x"fe"),
  1542 => (x"e8",x"c0",x"85",x"c2"),
  1543 => (x"80",x"c1",x"48",x"66"),
  1544 => (x"58",x"a6",x"ec",x"c0"),
  1545 => (x"49",x"66",x"ec",x"c0"),
  1546 => (x"a9",x"70",x"81",x"c1"),
  1547 => (x"87",x"c8",x"c0",x"02"),
  1548 => (x"c0",x"48",x"a6",x"d8"),
  1549 => (x"87",x"c5",x"c0",x"78"),
  1550 => (x"c1",x"48",x"a6",x"d8"),
  1551 => (x"1e",x"66",x"d8",x"78"),
  1552 => (x"c0",x"49",x"a4",x"c2"),
  1553 => (x"88",x"71",x"48",x"e0"),
  1554 => (x"75",x"1e",x"49",x"70"),
  1555 => (x"f9",x"db",x"ff",x"49"),
  1556 => (x"c0",x"86",x"c8",x"87"),
  1557 => (x"ff",x"01",x"a8",x"b7"),
  1558 => (x"e8",x"c0",x"87",x"c0"),
  1559 => (x"d1",x"c0",x"02",x"66"),
  1560 => (x"c9",x"49",x"6e",x"87"),
  1561 => (x"66",x"e8",x"c0",x"81"),
  1562 => (x"c1",x"48",x"6e",x"51"),
  1563 => (x"c0",x"78",x"df",x"cf"),
  1564 => (x"49",x"6e",x"87",x"cc"),
  1565 => (x"51",x"c2",x"81",x"c9"),
  1566 => (x"d0",x"c1",x"48",x"6e"),
  1567 => (x"7e",x"c1",x"78",x"d3"),
  1568 => (x"ff",x"87",x"c6",x"c0"),
  1569 => (x"70",x"87",x"ef",x"da"),
  1570 => (x"c0",x"02",x"6e",x"4c"),
  1571 => (x"66",x"c4",x"87",x"f5"),
  1572 => (x"a8",x"66",x"c8",x"48"),
  1573 => (x"87",x"cb",x"c0",x"04"),
  1574 => (x"c1",x"48",x"66",x"c4"),
  1575 => (x"58",x"a6",x"c8",x"80"),
  1576 => (x"c8",x"87",x"e0",x"c0"),
  1577 => (x"88",x"c1",x"48",x"66"),
  1578 => (x"c0",x"58",x"a6",x"cc"),
  1579 => (x"c6",x"c1",x"87",x"d5"),
  1580 => (x"c8",x"c0",x"05",x"ac"),
  1581 => (x"48",x"66",x"cc",x"87"),
  1582 => (x"a6",x"d0",x"80",x"c1"),
  1583 => (x"f5",x"d9",x"ff",x"58"),
  1584 => (x"d0",x"4c",x"70",x"87"),
  1585 => (x"80",x"c1",x"48",x"66"),
  1586 => (x"74",x"58",x"a6",x"d4"),
  1587 => (x"cb",x"c0",x"02",x"9c"),
  1588 => (x"48",x"66",x"c4",x"87"),
  1589 => (x"a8",x"66",x"c8",x"c1"),
  1590 => (x"87",x"ff",x"f2",x"04"),
  1591 => (x"87",x"cd",x"d9",x"ff"),
  1592 => (x"c7",x"48",x"66",x"c4"),
  1593 => (x"e5",x"c0",x"03",x"a8"),
  1594 => (x"cc",x"fd",x"c3",x"87"),
  1595 => (x"c4",x"78",x"c0",x"48"),
  1596 => (x"91",x"cb",x"49",x"66"),
  1597 => (x"81",x"66",x"c0",x"c1"),
  1598 => (x"6a",x"4a",x"a1",x"c4"),
  1599 => (x"79",x"52",x"c0",x"4a"),
  1600 => (x"c1",x"48",x"66",x"c4"),
  1601 => (x"58",x"a6",x"c8",x"80"),
  1602 => (x"ff",x"04",x"a8",x"c7"),
  1603 => (x"d0",x"ff",x"87",x"db"),
  1604 => (x"87",x"f5",x"e0",x"8e"),
  1605 => (x"1e",x"00",x"20",x"3a"),
  1606 => (x"4b",x"71",x"1e",x"73"),
  1607 => (x"87",x"c6",x"02",x"9b"),
  1608 => (x"48",x"c8",x"fd",x"c3"),
  1609 => (x"1e",x"c7",x"78",x"c0"),
  1610 => (x"bf",x"c8",x"fd",x"c3"),
  1611 => (x"e9",x"c1",x"1e",x"49"),
  1612 => (x"fd",x"c3",x"1e",x"d7"),
  1613 => (x"ee",x"49",x"bf",x"c4"),
  1614 => (x"86",x"cc",x"87",x"f4"),
  1615 => (x"bf",x"c4",x"fd",x"c3"),
  1616 => (x"87",x"f3",x"e9",x"49"),
  1617 => (x"c8",x"02",x"9b",x"73"),
  1618 => (x"d7",x"e9",x"c1",x"87"),
  1619 => (x"c2",x"e7",x"c0",x"49"),
  1620 => (x"f8",x"df",x"ff",x"87"),
  1621 => (x"1e",x"73",x"1e",x"87"),
  1622 => (x"4b",x"ff",x"c3",x"1e"),
  1623 => (x"fc",x"4a",x"d4",x"ff"),
  1624 => (x"98",x"c1",x"48",x"bf"),
  1625 => (x"02",x"6e",x"7e",x"70"),
  1626 => (x"ff",x"87",x"fb",x"c0"),
  1627 => (x"c1",x"c1",x"48",x"d0"),
  1628 => (x"7a",x"d2",x"c2",x"78"),
  1629 => (x"f0",x"c3",x"7a",x"73"),
  1630 => (x"ff",x"48",x"49",x"d3"),
  1631 => (x"73",x"50",x"6a",x"80"),
  1632 => (x"73",x"51",x"6a",x"7a"),
  1633 => (x"6a",x"80",x"c1",x"7a"),
  1634 => (x"6a",x"7a",x"73",x"50"),
  1635 => (x"6a",x"7a",x"73",x"50"),
  1636 => (x"6a",x"7a",x"73",x"49"),
  1637 => (x"6a",x"7a",x"73",x"50"),
  1638 => (x"dc",x"f0",x"c3",x"50"),
  1639 => (x"d0",x"ff",x"59",x"97"),
  1640 => (x"78",x"c0",x"c1",x"48"),
  1641 => (x"f0",x"c3",x"87",x"d7"),
  1642 => (x"ff",x"48",x"49",x"d3"),
  1643 => (x"51",x"50",x"c0",x"80"),
  1644 => (x"50",x"c0",x"80",x"c1"),
  1645 => (x"50",x"c1",x"50",x"d9"),
  1646 => (x"c3",x"50",x"e2",x"c0"),
  1647 => (x"d9",x"f0",x"c3",x"50"),
  1648 => (x"f8",x"50",x"c0",x"48"),
  1649 => (x"de",x"ff",x"26",x"80"),
  1650 => (x"c7",x"1e",x"87",x"c3"),
  1651 => (x"49",x"c1",x"87",x"cb"),
  1652 => (x"fe",x"87",x"c4",x"fd"),
  1653 => (x"70",x"87",x"d4",x"e6"),
  1654 => (x"87",x"cd",x"02",x"98"),
  1655 => (x"87",x"d1",x"ef",x"fe"),
  1656 => (x"c4",x"02",x"98",x"70"),
  1657 => (x"c2",x"4a",x"c1",x"87"),
  1658 => (x"72",x"4a",x"c0",x"87"),
  1659 => (x"87",x"ce",x"05",x"9a"),
  1660 => (x"e8",x"c1",x"1e",x"c0"),
  1661 => (x"f0",x"c0",x"49",x"db"),
  1662 => (x"86",x"c4",x"87",x"f4"),
  1663 => (x"1e",x"c0",x"87",x"fe"),
  1664 => (x"49",x"e6",x"e8",x"c1"),
  1665 => (x"87",x"e6",x"f0",x"c0"),
  1666 => (x"fb",x"c1",x"1e",x"c0"),
  1667 => (x"49",x"70",x"87",x"c6"),
  1668 => (x"87",x"da",x"f0",x"c0"),
  1669 => (x"f8",x"87",x"c1",x"c3"),
  1670 => (x"53",x"4f",x"26",x"8e"),
  1671 => (x"61",x"66",x"20",x"44"),
  1672 => (x"64",x"65",x"6c",x"69"),
  1673 => (x"6f",x"42",x"00",x"2e"),
  1674 => (x"6e",x"69",x"74",x"6f"),
  1675 => (x"2e",x"2e",x"2e",x"67"),
  1676 => (x"fd",x"c3",x"1e",x"00"),
  1677 => (x"78",x"c0",x"48",x"c8"),
  1678 => (x"48",x"c4",x"fd",x"c3"),
  1679 => (x"c9",x"fe",x"78",x"c0"),
  1680 => (x"f6",x"fd",x"c1",x"87"),
  1681 => (x"26",x"48",x"c0",x"87"),
  1682 => (x"45",x"20",x"80",x"4f"),
  1683 => (x"00",x"74",x"69",x"78"),
  1684 => (x"61",x"42",x"20",x"80"),
  1685 => (x"8f",x"00",x"6b",x"63"),
  1686 => (x"5d",x"00",x"00",x"13"),
  1687 => (x"00",x"00",x"00",x"3f"),
  1688 => (x"13",x"8f",x"00",x"00"),
  1689 => (x"3f",x"7b",x"00",x"00"),
  1690 => (x"00",x"00",x"00",x"00"),
  1691 => (x"00",x"13",x"8f",x"00"),
  1692 => (x"00",x"3f",x"99",x"00"),
  1693 => (x"00",x"00",x"00",x"00"),
  1694 => (x"00",x"00",x"13",x"8f"),
  1695 => (x"00",x"00",x"3f",x"b7"),
  1696 => (x"8f",x"00",x"00",x"00"),
  1697 => (x"d5",x"00",x"00",x"13"),
  1698 => (x"00",x"00",x"00",x"3f"),
  1699 => (x"13",x"8f",x"00",x"00"),
  1700 => (x"3f",x"f3",x"00",x"00"),
  1701 => (x"00",x"00",x"00",x"00"),
  1702 => (x"00",x"13",x"8f",x"00"),
  1703 => (x"00",x"40",x"11",x"00"),
  1704 => (x"00",x"00",x"00",x"00"),
  1705 => (x"00",x"00",x"13",x"8f"),
  1706 => (x"00",x"00",x"00",x"00"),
  1707 => (x"2a",x"00",x"00",x"00"),
  1708 => (x"00",x"00",x"00",x"14"),
  1709 => (x"00",x"00",x"00",x"00"),
  1710 => (x"6f",x"4c",x"00",x"00"),
  1711 => (x"2a",x"20",x"64",x"61"),
  1712 => (x"fe",x"1e",x"00",x"2e"),
  1713 => (x"78",x"c0",x"48",x"f0"),
  1714 => (x"09",x"79",x"09",x"cd"),
  1715 => (x"1e",x"1e",x"4f",x"26"),
  1716 => (x"7e",x"bf",x"f0",x"fe"),
  1717 => (x"4f",x"26",x"26",x"48"),
  1718 => (x"48",x"f0",x"fe",x"1e"),
  1719 => (x"4f",x"26",x"78",x"c1"),
  1720 => (x"48",x"f0",x"fe",x"1e"),
  1721 => (x"4f",x"26",x"78",x"c0"),
  1722 => (x"c0",x"4a",x"71",x"1e"),
  1723 => (x"4f",x"26",x"52",x"52"),
  1724 => (x"5c",x"5b",x"5e",x"0e"),
  1725 => (x"86",x"f4",x"0e",x"5d"),
  1726 => (x"6d",x"97",x"4d",x"71"),
  1727 => (x"4c",x"a5",x"c1",x"7e"),
  1728 => (x"c8",x"48",x"6c",x"97"),
  1729 => (x"48",x"6e",x"58",x"a6"),
  1730 => (x"05",x"a8",x"66",x"c4"),
  1731 => (x"48",x"ff",x"87",x"c5"),
  1732 => (x"ff",x"87",x"e6",x"c0"),
  1733 => (x"a5",x"c2",x"87",x"ca"),
  1734 => (x"4b",x"6c",x"97",x"49"),
  1735 => (x"97",x"4b",x"a3",x"71"),
  1736 => (x"6c",x"97",x"4b",x"6b"),
  1737 => (x"c1",x"48",x"6e",x"7e"),
  1738 => (x"58",x"a6",x"c8",x"80"),
  1739 => (x"a6",x"cc",x"98",x"c7"),
  1740 => (x"7c",x"97",x"70",x"58"),
  1741 => (x"73",x"87",x"e1",x"fe"),
  1742 => (x"26",x"8e",x"f4",x"48"),
  1743 => (x"26",x"4c",x"26",x"4d"),
  1744 => (x"0e",x"4f",x"26",x"4b"),
  1745 => (x"0e",x"5c",x"5b",x"5e"),
  1746 => (x"4c",x"71",x"86",x"f4"),
  1747 => (x"c3",x"4a",x"66",x"d8"),
  1748 => (x"a4",x"c2",x"9a",x"ff"),
  1749 => (x"49",x"6c",x"97",x"4b"),
  1750 => (x"72",x"49",x"a1",x"73"),
  1751 => (x"7e",x"6c",x"97",x"51"),
  1752 => (x"80",x"c1",x"48",x"6e"),
  1753 => (x"c7",x"58",x"a6",x"c8"),
  1754 => (x"58",x"a6",x"cc",x"98"),
  1755 => (x"8e",x"f4",x"54",x"70"),
  1756 => (x"1e",x"87",x"ca",x"ff"),
  1757 => (x"87",x"e8",x"fd",x"1e"),
  1758 => (x"49",x"4a",x"bf",x"e0"),
  1759 => (x"99",x"c0",x"e0",x"c0"),
  1760 => (x"72",x"87",x"cb",x"02"),
  1761 => (x"ef",x"c0",x"c4",x"1e"),
  1762 => (x"87",x"f7",x"fe",x"49"),
  1763 => (x"fd",x"fc",x"86",x"c4"),
  1764 => (x"fd",x"7e",x"70",x"87"),
  1765 => (x"26",x"26",x"87",x"c2"),
  1766 => (x"c0",x"c4",x"1e",x"4f"),
  1767 => (x"c7",x"fd",x"49",x"ef"),
  1768 => (x"f3",x"ed",x"c1",x"87"),
  1769 => (x"87",x"da",x"fc",x"49"),
  1770 => (x"26",x"87",x"f8",x"c4"),
  1771 => (x"5b",x"5e",x"0e",x"4f"),
  1772 => (x"c4",x"0e",x"5d",x"5c"),
  1773 => (x"4a",x"bf",x"ce",x"c1"),
  1774 => (x"bf",x"c1",x"f0",x"c1"),
  1775 => (x"bc",x"72",x"4c",x"49"),
  1776 => (x"db",x"fc",x"4d",x"71"),
  1777 => (x"74",x"4b",x"c0",x"87"),
  1778 => (x"02",x"99",x"d0",x"49"),
  1779 => (x"49",x"75",x"87",x"d5"),
  1780 => (x"1e",x"71",x"99",x"d0"),
  1781 => (x"f5",x"c1",x"1e",x"c0"),
  1782 => (x"82",x"73",x"4a",x"f2"),
  1783 => (x"e4",x"c0",x"49",x"12"),
  1784 => (x"c1",x"86",x"c8",x"87"),
  1785 => (x"c8",x"83",x"2d",x"2c"),
  1786 => (x"da",x"ff",x"04",x"ab"),
  1787 => (x"87",x"e8",x"fb",x"87"),
  1788 => (x"48",x"c1",x"f0",x"c1"),
  1789 => (x"bf",x"ce",x"c1",x"c4"),
  1790 => (x"26",x"4d",x"26",x"78"),
  1791 => (x"26",x"4b",x"26",x"4c"),
  1792 => (x"00",x"00",x"00",x"4f"),
  1793 => (x"d0",x"ff",x"1e",x"00"),
  1794 => (x"78",x"e1",x"c8",x"48"),
  1795 => (x"c5",x"48",x"d4",x"ff"),
  1796 => (x"02",x"66",x"c4",x"78"),
  1797 => (x"e0",x"c3",x"87",x"c3"),
  1798 => (x"02",x"66",x"c8",x"78"),
  1799 => (x"d4",x"ff",x"87",x"c6"),
  1800 => (x"78",x"f0",x"c3",x"48"),
  1801 => (x"71",x"48",x"d4",x"ff"),
  1802 => (x"48",x"d0",x"ff",x"78"),
  1803 => (x"c0",x"78",x"e1",x"c8"),
  1804 => (x"4f",x"26",x"78",x"e0"),
  1805 => (x"c4",x"1e",x"73",x"1e"),
  1806 => (x"fa",x"49",x"ef",x"c0"),
  1807 => (x"4a",x"70",x"87",x"f2"),
  1808 => (x"04",x"aa",x"b7",x"c0"),
  1809 => (x"c3",x"87",x"cf",x"c2"),
  1810 => (x"c9",x"05",x"aa",x"e0"),
  1811 => (x"df",x"f3",x"c1",x"87"),
  1812 => (x"c2",x"78",x"c1",x"48"),
  1813 => (x"49",x"72",x"87",x"c0"),
  1814 => (x"02",x"99",x"c0",x"c2"),
  1815 => (x"f3",x"c1",x"87",x"c9"),
  1816 => (x"78",x"c1",x"48",x"db"),
  1817 => (x"c1",x"9a",x"ff",x"fd"),
  1818 => (x"02",x"bf",x"df",x"f3"),
  1819 => (x"4b",x"72",x"87",x"c7"),
  1820 => (x"c2",x"b3",x"c0",x"c2"),
  1821 => (x"c1",x"4b",x"72",x"87"),
  1822 => (x"02",x"bf",x"db",x"f3"),
  1823 => (x"73",x"87",x"e0",x"c0"),
  1824 => (x"29",x"b7",x"c4",x"49"),
  1825 => (x"f2",x"f4",x"c1",x"91"),
  1826 => (x"cf",x"4a",x"73",x"81"),
  1827 => (x"c1",x"92",x"c2",x"9a"),
  1828 => (x"70",x"30",x"72",x"48"),
  1829 => (x"72",x"ba",x"ff",x"4a"),
  1830 => (x"70",x"98",x"69",x"48"),
  1831 => (x"73",x"87",x"db",x"79"),
  1832 => (x"29",x"b7",x"c4",x"49"),
  1833 => (x"f2",x"f4",x"c1",x"91"),
  1834 => (x"cf",x"4a",x"73",x"81"),
  1835 => (x"c3",x"92",x"c2",x"9a"),
  1836 => (x"70",x"30",x"72",x"48"),
  1837 => (x"b0",x"69",x"48",x"4a"),
  1838 => (x"f3",x"c1",x"79",x"70"),
  1839 => (x"78",x"c0",x"48",x"df"),
  1840 => (x"48",x"db",x"f3",x"c1"),
  1841 => (x"c0",x"c4",x"78",x"c0"),
  1842 => (x"e3",x"f8",x"49",x"ef"),
  1843 => (x"c0",x"4a",x"70",x"87"),
  1844 => (x"fd",x"03",x"aa",x"b7"),
  1845 => (x"48",x"c0",x"87",x"f1"),
  1846 => (x"00",x"87",x"e2",x"fc"),
  1847 => (x"00",x"00",x"00",x"00"),
  1848 => (x"1e",x"00",x"00",x"00"),
  1849 => (x"49",x"72",x"4a",x"c0"),
  1850 => (x"f4",x"c1",x"91",x"c4"),
  1851 => (x"79",x"c0",x"81",x"f2"),
  1852 => (x"b7",x"d0",x"82",x"c1"),
  1853 => (x"87",x"ee",x"04",x"aa"),
  1854 => (x"5e",x"0e",x"4f",x"26"),
  1855 => (x"0e",x"5d",x"5c",x"5b"),
  1856 => (x"db",x"f7",x"4d",x"71"),
  1857 => (x"c4",x"4a",x"75",x"87"),
  1858 => (x"c1",x"92",x"2a",x"b7"),
  1859 => (x"75",x"82",x"f2",x"f4"),
  1860 => (x"c2",x"9c",x"cf",x"4c"),
  1861 => (x"4b",x"49",x"6a",x"94"),
  1862 => (x"9b",x"c3",x"2b",x"74"),
  1863 => (x"30",x"74",x"48",x"c2"),
  1864 => (x"bc",x"ff",x"4c",x"70"),
  1865 => (x"98",x"71",x"48",x"74"),
  1866 => (x"eb",x"f6",x"7a",x"70"),
  1867 => (x"fb",x"48",x"73",x"87"),
  1868 => (x"00",x"00",x"87",x"c7"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"00",x"00"),
  1871 => (x"00",x"00",x"00",x"00"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"00",x"00"),
  1875 => (x"00",x"00",x"00",x"00"),
  1876 => (x"00",x"00",x"00",x"00"),
  1877 => (x"00",x"00",x"00",x"00"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"00",x"00",x"00",x"00"),
  1883 => (x"00",x"00",x"00",x"00"),
  1884 => (x"1e",x"16",x"00",x"00"),
  1885 => (x"36",x"2e",x"25",x"26"),
  1886 => (x"ff",x"1e",x"3e",x"3d"),
  1887 => (x"e1",x"c8",x"48",x"d0"),
  1888 => (x"ff",x"48",x"71",x"78"),
  1889 => (x"26",x"78",x"08",x"d4"),
  1890 => (x"d0",x"ff",x"1e",x"4f"),
  1891 => (x"78",x"e1",x"c8",x"48"),
  1892 => (x"d4",x"ff",x"48",x"71"),
  1893 => (x"66",x"c4",x"78",x"08"),
  1894 => (x"08",x"d4",x"ff",x"48"),
  1895 => (x"1e",x"4f",x"26",x"78"),
  1896 => (x"66",x"c4",x"4a",x"71"),
  1897 => (x"49",x"72",x"1e",x"49"),
  1898 => (x"ff",x"87",x"de",x"ff"),
  1899 => (x"e0",x"c0",x"48",x"d0"),
  1900 => (x"4f",x"26",x"26",x"78"),
  1901 => (x"c4",x"4a",x"71",x"1e"),
  1902 => (x"e0",x"c1",x"1e",x"66"),
  1903 => (x"c8",x"ff",x"49",x"a2"),
  1904 => (x"49",x"66",x"c8",x"87"),
  1905 => (x"ff",x"29",x"b7",x"c8"),
  1906 => (x"78",x"71",x"48",x"d4"),
  1907 => (x"c0",x"48",x"d0",x"ff"),
  1908 => (x"26",x"26",x"78",x"e0"),
  1909 => (x"1e",x"73",x"1e",x"4f"),
  1910 => (x"e2",x"c0",x"4b",x"71"),
  1911 => (x"87",x"da",x"fe",x"49"),
  1912 => (x"48",x"13",x"4a",x"c7"),
  1913 => (x"78",x"08",x"d4",x"ff"),
  1914 => (x"8a",x"c1",x"49",x"72"),
  1915 => (x"f1",x"05",x"99",x"71"),
  1916 => (x"48",x"d0",x"ff",x"87"),
  1917 => (x"c4",x"78",x"e0",x"c0"),
  1918 => (x"26",x"4d",x"26",x"87"),
  1919 => (x"26",x"4b",x"26",x"4c"),
  1920 => (x"d4",x"ff",x"1e",x"4f"),
  1921 => (x"7a",x"ff",x"c3",x"4a"),
  1922 => (x"c8",x"48",x"d0",x"ff"),
  1923 => (x"7a",x"de",x"78",x"e1"),
  1924 => (x"bf",x"f9",x"c0",x"c4"),
  1925 => (x"c8",x"48",x"49",x"7a"),
  1926 => (x"71",x"7a",x"70",x"28"),
  1927 => (x"70",x"28",x"d0",x"48"),
  1928 => (x"d8",x"48",x"71",x"7a"),
  1929 => (x"ff",x"7a",x"70",x"28"),
  1930 => (x"e0",x"c0",x"48",x"d0"),
  1931 => (x"0e",x"4f",x"26",x"78"),
  1932 => (x"5d",x"5c",x"5b",x"5e"),
  1933 => (x"c4",x"4c",x"71",x"0e"),
  1934 => (x"4d",x"bf",x"f9",x"c0"),
  1935 => (x"d0",x"2b",x"74",x"4b"),
  1936 => (x"83",x"c1",x"9b",x"66"),
  1937 => (x"04",x"ab",x"66",x"d4"),
  1938 => (x"4b",x"c0",x"87",x"c2"),
  1939 => (x"66",x"d0",x"4a",x"74"),
  1940 => (x"ff",x"31",x"72",x"49"),
  1941 => (x"73",x"99",x"75",x"b9"),
  1942 => (x"70",x"30",x"72",x"48"),
  1943 => (x"b0",x"71",x"48",x"4a"),
  1944 => (x"58",x"fd",x"c0",x"c4"),
  1945 => (x"26",x"87",x"da",x"fe"),
  1946 => (x"26",x"4c",x"26",x"4d"),
  1947 => (x"1e",x"4f",x"26",x"4b"),
  1948 => (x"c8",x"48",x"d0",x"ff"),
  1949 => (x"48",x"71",x"78",x"c9"),
  1950 => (x"78",x"08",x"d4",x"ff"),
  1951 => (x"71",x"1e",x"4f",x"26"),
  1952 => (x"87",x"eb",x"49",x"4a"),
  1953 => (x"c8",x"48",x"d0",x"ff"),
  1954 => (x"1e",x"4f",x"26",x"78"),
  1955 => (x"4b",x"71",x"1e",x"73"),
  1956 => (x"bf",x"c9",x"c1",x"c4"),
  1957 => (x"c2",x"87",x"c3",x"02"),
  1958 => (x"d0",x"ff",x"87",x"eb"),
  1959 => (x"78",x"c9",x"c8",x"48"),
  1960 => (x"e0",x"c0",x"49",x"73"),
  1961 => (x"48",x"d4",x"ff",x"b1"),
  1962 => (x"c0",x"c4",x"78",x"71"),
  1963 => (x"78",x"c0",x"48",x"fd"),
  1964 => (x"c5",x"02",x"66",x"c8"),
  1965 => (x"49",x"ff",x"c3",x"87"),
  1966 => (x"49",x"c0",x"87",x"c2"),
  1967 => (x"59",x"c5",x"c1",x"c4"),
  1968 => (x"c6",x"02",x"66",x"cc"),
  1969 => (x"d5",x"d5",x"c5",x"87"),
  1970 => (x"cf",x"87",x"c4",x"4a"),
  1971 => (x"c4",x"4a",x"ff",x"ff"),
  1972 => (x"c4",x"5a",x"c9",x"c1"),
  1973 => (x"c1",x"48",x"c9",x"c1"),
  1974 => (x"26",x"87",x"c4",x"78"),
  1975 => (x"26",x"4c",x"26",x"4d"),
  1976 => (x"0e",x"4f",x"26",x"4b"),
  1977 => (x"5d",x"5c",x"5b",x"5e"),
  1978 => (x"c4",x"4a",x"71",x"0e"),
  1979 => (x"4c",x"bf",x"c5",x"c1"),
  1980 => (x"cb",x"02",x"9a",x"72"),
  1981 => (x"91",x"c8",x"49",x"87"),
  1982 => (x"4b",x"c1",x"fa",x"c1"),
  1983 => (x"87",x"c4",x"83",x"71"),
  1984 => (x"4b",x"c1",x"fe",x"c1"),
  1985 => (x"49",x"13",x"4d",x"c0"),
  1986 => (x"c1",x"c4",x"99",x"74"),
  1987 => (x"ff",x"b9",x"bf",x"c1"),
  1988 => (x"78",x"71",x"48",x"d4"),
  1989 => (x"85",x"2c",x"b7",x"c1"),
  1990 => (x"04",x"ad",x"b7",x"c8"),
  1991 => (x"c0",x"c4",x"87",x"e8"),
  1992 => (x"c8",x"48",x"bf",x"fd"),
  1993 => (x"c1",x"c1",x"c4",x"80"),
  1994 => (x"87",x"ef",x"fe",x"58"),
  1995 => (x"71",x"1e",x"73",x"1e"),
  1996 => (x"9a",x"4a",x"13",x"4b"),
  1997 => (x"72",x"87",x"cb",x"02"),
  1998 => (x"87",x"e7",x"fe",x"49"),
  1999 => (x"05",x"9a",x"4a",x"13"),
  2000 => (x"da",x"fe",x"87",x"f5"),
  2001 => (x"c0",x"c4",x"1e",x"87"),
  2002 => (x"c4",x"49",x"bf",x"fd"),
  2003 => (x"c1",x"48",x"fd",x"c0"),
  2004 => (x"c0",x"c4",x"78",x"a1"),
  2005 => (x"db",x"03",x"a9",x"b7"),
  2006 => (x"48",x"d4",x"ff",x"87"),
  2007 => (x"bf",x"c1",x"c1",x"c4"),
  2008 => (x"fd",x"c0",x"c4",x"78"),
  2009 => (x"c0",x"c4",x"49",x"bf"),
  2010 => (x"a1",x"c1",x"48",x"fd"),
  2011 => (x"b7",x"c0",x"c4",x"78"),
  2012 => (x"87",x"e5",x"04",x"a9"),
  2013 => (x"c8",x"48",x"d0",x"ff"),
  2014 => (x"c9",x"c1",x"c4",x"78"),
  2015 => (x"26",x"78",x"c0",x"48"),
  2016 => (x"00",x"00",x"00",x"4f"),
  2017 => (x"00",x"00",x"00",x"00"),
  2018 => (x"00",x"00",x"00",x"00"),
  2019 => (x"00",x"00",x"5f",x"5f"),
  2020 => (x"03",x"03",x"00",x"00"),
  2021 => (x"00",x"03",x"03",x"00"),
  2022 => (x"7f",x"7f",x"14",x"00"),
  2023 => (x"14",x"7f",x"7f",x"14"),
  2024 => (x"2e",x"24",x"00",x"00"),
  2025 => (x"12",x"3a",x"6b",x"6b"),
  2026 => (x"36",x"6a",x"4c",x"00"),
  2027 => (x"32",x"56",x"6c",x"18"),
  2028 => (x"4f",x"7e",x"30",x"00"),
  2029 => (x"68",x"3a",x"77",x"59"),
  2030 => (x"04",x"00",x"00",x"40"),
  2031 => (x"00",x"00",x"03",x"07"),
  2032 => (x"1c",x"00",x"00",x"00"),
  2033 => (x"00",x"41",x"63",x"3e"),
  2034 => (x"41",x"00",x"00",x"00"),
  2035 => (x"00",x"1c",x"3e",x"63"),
  2036 => (x"3e",x"2a",x"08",x"00"),
  2037 => (x"2a",x"3e",x"1c",x"1c"),
  2038 => (x"08",x"08",x"00",x"08"),
  2039 => (x"08",x"08",x"3e",x"3e"),
  2040 => (x"80",x"00",x"00",x"00"),
  2041 => (x"00",x"00",x"60",x"e0"),
  2042 => (x"08",x"08",x"00",x"00"),
  2043 => (x"08",x"08",x"08",x"08"),
  2044 => (x"00",x"00",x"00",x"00"),
  2045 => (x"00",x"00",x"60",x"60"),
  2046 => (x"30",x"60",x"40",x"00"),
  2047 => (x"03",x"06",x"0c",x"18"),
  2048 => (x"7f",x"3e",x"00",x"01"),
  2049 => (x"3e",x"7f",x"4d",x"59"),
  2050 => (x"06",x"04",x"00",x"00"),
  2051 => (x"00",x"00",x"7f",x"7f"),
  2052 => (x"63",x"42",x"00",x"00"),
  2053 => (x"46",x"4f",x"59",x"71"),
  2054 => (x"63",x"22",x"00",x"00"),
  2055 => (x"36",x"7f",x"49",x"49"),
  2056 => (x"16",x"1c",x"18",x"00"),
  2057 => (x"10",x"7f",x"7f",x"13"),
  2058 => (x"67",x"27",x"00",x"00"),
  2059 => (x"39",x"7d",x"45",x"45"),
  2060 => (x"7e",x"3c",x"00",x"00"),
  2061 => (x"30",x"79",x"49",x"4b"),
  2062 => (x"01",x"01",x"00",x"00"),
  2063 => (x"07",x"0f",x"79",x"71"),
  2064 => (x"7f",x"36",x"00",x"00"),
  2065 => (x"36",x"7f",x"49",x"49"),
  2066 => (x"4f",x"06",x"00",x"00"),
  2067 => (x"1e",x"3f",x"69",x"49"),
  2068 => (x"00",x"00",x"00",x"00"),
  2069 => (x"00",x"00",x"66",x"66"),
  2070 => (x"80",x"00",x"00",x"00"),
  2071 => (x"00",x"00",x"66",x"e6"),
  2072 => (x"08",x"08",x"00",x"00"),
  2073 => (x"22",x"22",x"14",x"14"),
  2074 => (x"14",x"14",x"00",x"00"),
  2075 => (x"14",x"14",x"14",x"14"),
  2076 => (x"22",x"22",x"00",x"00"),
  2077 => (x"08",x"08",x"14",x"14"),
  2078 => (x"03",x"02",x"00",x"00"),
  2079 => (x"06",x"0f",x"59",x"51"),
  2080 => (x"41",x"7f",x"3e",x"00"),
  2081 => (x"1e",x"1f",x"55",x"5d"),
  2082 => (x"7f",x"7e",x"00",x"00"),
  2083 => (x"7e",x"7f",x"09",x"09"),
  2084 => (x"7f",x"7f",x"00",x"00"),
  2085 => (x"36",x"7f",x"49",x"49"),
  2086 => (x"3e",x"1c",x"00",x"00"),
  2087 => (x"41",x"41",x"41",x"63"),
  2088 => (x"7f",x"7f",x"00",x"00"),
  2089 => (x"1c",x"3e",x"63",x"41"),
  2090 => (x"7f",x"7f",x"00",x"00"),
  2091 => (x"41",x"41",x"49",x"49"),
  2092 => (x"7f",x"7f",x"00",x"00"),
  2093 => (x"01",x"01",x"09",x"09"),
  2094 => (x"7f",x"3e",x"00",x"00"),
  2095 => (x"7a",x"7b",x"49",x"41"),
  2096 => (x"7f",x"7f",x"00",x"00"),
  2097 => (x"7f",x"7f",x"08",x"08"),
  2098 => (x"41",x"00",x"00",x"00"),
  2099 => (x"00",x"41",x"7f",x"7f"),
  2100 => (x"60",x"20",x"00",x"00"),
  2101 => (x"3f",x"7f",x"40",x"40"),
  2102 => (x"08",x"7f",x"7f",x"00"),
  2103 => (x"41",x"63",x"36",x"1c"),
  2104 => (x"7f",x"7f",x"00",x"00"),
  2105 => (x"40",x"40",x"40",x"40"),
  2106 => (x"06",x"7f",x"7f",x"00"),
  2107 => (x"7f",x"7f",x"06",x"0c"),
  2108 => (x"06",x"7f",x"7f",x"00"),
  2109 => (x"7f",x"7f",x"18",x"0c"),
  2110 => (x"7f",x"3e",x"00",x"00"),
  2111 => (x"3e",x"7f",x"41",x"41"),
  2112 => (x"7f",x"7f",x"00",x"00"),
  2113 => (x"06",x"0f",x"09",x"09"),
  2114 => (x"41",x"7f",x"3e",x"00"),
  2115 => (x"40",x"7e",x"7f",x"61"),
  2116 => (x"7f",x"7f",x"00",x"00"),
  2117 => (x"66",x"7f",x"19",x"09"),
  2118 => (x"6f",x"26",x"00",x"00"),
  2119 => (x"32",x"7b",x"59",x"4d"),
  2120 => (x"01",x"01",x"00",x"00"),
  2121 => (x"01",x"01",x"7f",x"7f"),
  2122 => (x"7f",x"3f",x"00",x"00"),
  2123 => (x"3f",x"7f",x"40",x"40"),
  2124 => (x"3f",x"0f",x"00",x"00"),
  2125 => (x"0f",x"3f",x"70",x"70"),
  2126 => (x"30",x"7f",x"7f",x"00"),
  2127 => (x"7f",x"7f",x"30",x"18"),
  2128 => (x"36",x"63",x"41",x"00"),
  2129 => (x"63",x"36",x"1c",x"1c"),
  2130 => (x"06",x"03",x"01",x"41"),
  2131 => (x"03",x"06",x"7c",x"7c"),
  2132 => (x"59",x"71",x"61",x"01"),
  2133 => (x"41",x"43",x"47",x"4d"),
  2134 => (x"7f",x"00",x"00",x"00"),
  2135 => (x"00",x"41",x"41",x"7f"),
  2136 => (x"06",x"03",x"01",x"00"),
  2137 => (x"60",x"30",x"18",x"0c"),
  2138 => (x"41",x"00",x"00",x"40"),
  2139 => (x"00",x"7f",x"7f",x"41"),
  2140 => (x"06",x"0c",x"08",x"00"),
  2141 => (x"08",x"0c",x"06",x"03"),
  2142 => (x"80",x"80",x"80",x"00"),
  2143 => (x"80",x"80",x"80",x"80"),
  2144 => (x"00",x"00",x"00",x"00"),
  2145 => (x"00",x"04",x"07",x"03"),
  2146 => (x"74",x"20",x"00",x"00"),
  2147 => (x"78",x"7c",x"54",x"54"),
  2148 => (x"7f",x"7f",x"00",x"00"),
  2149 => (x"38",x"7c",x"44",x"44"),
  2150 => (x"7c",x"38",x"00",x"00"),
  2151 => (x"00",x"44",x"44",x"44"),
  2152 => (x"7c",x"38",x"00",x"00"),
  2153 => (x"7f",x"7f",x"44",x"44"),
  2154 => (x"7c",x"38",x"00",x"00"),
  2155 => (x"18",x"5c",x"54",x"54"),
  2156 => (x"7e",x"04",x"00",x"00"),
  2157 => (x"00",x"05",x"05",x"7f"),
  2158 => (x"bc",x"18",x"00",x"00"),
  2159 => (x"7c",x"fc",x"a4",x"a4"),
  2160 => (x"7f",x"7f",x"00",x"00"),
  2161 => (x"78",x"7c",x"04",x"04"),
  2162 => (x"00",x"00",x"00",x"00"),
  2163 => (x"00",x"40",x"7d",x"3d"),
  2164 => (x"80",x"80",x"00",x"00"),
  2165 => (x"00",x"7d",x"fd",x"80"),
  2166 => (x"7f",x"7f",x"00",x"00"),
  2167 => (x"44",x"6c",x"38",x"10"),
  2168 => (x"00",x"00",x"00",x"00"),
  2169 => (x"00",x"40",x"7f",x"3f"),
  2170 => (x"0c",x"7c",x"7c",x"00"),
  2171 => (x"78",x"7c",x"0c",x"18"),
  2172 => (x"7c",x"7c",x"00",x"00"),
  2173 => (x"78",x"7c",x"04",x"04"),
  2174 => (x"7c",x"38",x"00",x"00"),
  2175 => (x"38",x"7c",x"44",x"44"),
  2176 => (x"fc",x"fc",x"00",x"00"),
  2177 => (x"18",x"3c",x"24",x"24"),
  2178 => (x"3c",x"18",x"00",x"00"),
  2179 => (x"fc",x"fc",x"24",x"24"),
  2180 => (x"7c",x"7c",x"00",x"00"),
  2181 => (x"08",x"0c",x"04",x"04"),
  2182 => (x"5c",x"48",x"00",x"00"),
  2183 => (x"20",x"74",x"54",x"54"),
  2184 => (x"3f",x"04",x"00",x"00"),
  2185 => (x"00",x"44",x"44",x"7f"),
  2186 => (x"7c",x"3c",x"00",x"00"),
  2187 => (x"7c",x"7c",x"40",x"40"),
  2188 => (x"3c",x"1c",x"00",x"00"),
  2189 => (x"1c",x"3c",x"60",x"60"),
  2190 => (x"60",x"7c",x"3c",x"00"),
  2191 => (x"3c",x"7c",x"60",x"30"),
  2192 => (x"38",x"6c",x"44",x"00"),
  2193 => (x"44",x"6c",x"38",x"10"),
  2194 => (x"bc",x"1c",x"00",x"00"),
  2195 => (x"1c",x"3c",x"60",x"e0"),
  2196 => (x"64",x"44",x"00",x"00"),
  2197 => (x"44",x"4c",x"5c",x"74"),
  2198 => (x"08",x"08",x"00",x"00"),
  2199 => (x"41",x"41",x"77",x"3e"),
  2200 => (x"00",x"00",x"00",x"00"),
  2201 => (x"00",x"00",x"7f",x"7f"),
  2202 => (x"41",x"41",x"00",x"00"),
  2203 => (x"08",x"08",x"3e",x"77"),
  2204 => (x"01",x"01",x"02",x"00"),
  2205 => (x"01",x"02",x"02",x"03"),
  2206 => (x"7f",x"7f",x"7f",x"00"),
  2207 => (x"7f",x"7f",x"7f",x"7f"),
  2208 => (x"1c",x"08",x"08",x"00"),
  2209 => (x"7f",x"3e",x"3e",x"1c"),
  2210 => (x"3e",x"7f",x"7f",x"7f"),
  2211 => (x"08",x"1c",x"1c",x"3e"),
  2212 => (x"18",x"10",x"00",x"08"),
  2213 => (x"10",x"18",x"7c",x"7c"),
  2214 => (x"30",x"10",x"00",x"00"),
  2215 => (x"10",x"30",x"7c",x"7c"),
  2216 => (x"60",x"30",x"10",x"00"),
  2217 => (x"06",x"1e",x"78",x"60"),
  2218 => (x"3c",x"66",x"42",x"00"),
  2219 => (x"42",x"66",x"3c",x"18"),
  2220 => (x"6a",x"38",x"78",x"00"),
  2221 => (x"38",x"6c",x"c6",x"c2"),
  2222 => (x"00",x"00",x"60",x"00"),
  2223 => (x"60",x"00",x"00",x"60"),
  2224 => (x"5b",x"5e",x"0e",x"00"),
  2225 => (x"1e",x"0e",x"5d",x"5c"),
  2226 => (x"c1",x"c4",x"4c",x"71"),
  2227 => (x"c0",x"4d",x"bf",x"da"),
  2228 => (x"74",x"1e",x"c0",x"4b"),
  2229 => (x"87",x"c7",x"02",x"ab"),
  2230 => (x"c0",x"48",x"a6",x"c4"),
  2231 => (x"c4",x"87",x"c5",x"78"),
  2232 => (x"78",x"c1",x"48",x"a6"),
  2233 => (x"73",x"1e",x"66",x"c4"),
  2234 => (x"87",x"df",x"ee",x"49"),
  2235 => (x"e0",x"c0",x"86",x"c8"),
  2236 => (x"87",x"ef",x"ef",x"49"),
  2237 => (x"6a",x"4a",x"a5",x"c4"),
  2238 => (x"87",x"f0",x"f0",x"49"),
  2239 => (x"cb",x"87",x"c6",x"f1"),
  2240 => (x"c8",x"83",x"c1",x"85"),
  2241 => (x"ff",x"04",x"ab",x"b7"),
  2242 => (x"26",x"26",x"87",x"c7"),
  2243 => (x"26",x"4c",x"26",x"4d"),
  2244 => (x"1e",x"4f",x"26",x"4b"),
  2245 => (x"c1",x"c4",x"4a",x"71"),
  2246 => (x"c1",x"c4",x"5a",x"de"),
  2247 => (x"78",x"c7",x"48",x"de"),
  2248 => (x"87",x"dd",x"fe",x"49"),
  2249 => (x"73",x"1e",x"4f",x"26"),
  2250 => (x"c0",x"4a",x"71",x"1e"),
  2251 => (x"d3",x"03",x"aa",x"b7"),
  2252 => (x"c3",x"da",x"c2",x"87"),
  2253 => (x"87",x"c4",x"05",x"bf"),
  2254 => (x"87",x"c2",x"4b",x"c1"),
  2255 => (x"da",x"c2",x"4b",x"c0"),
  2256 => (x"87",x"c4",x"5b",x"c7"),
  2257 => (x"5a",x"c7",x"da",x"c2"),
  2258 => (x"bf",x"c3",x"da",x"c2"),
  2259 => (x"c1",x"9a",x"c1",x"4a"),
  2260 => (x"ec",x"49",x"a2",x"c0"),
  2261 => (x"48",x"fc",x"87",x"e8"),
  2262 => (x"bf",x"c3",x"da",x"c2"),
  2263 => (x"87",x"ef",x"fe",x"78"),
  2264 => (x"c3",x"da",x"c2",x"1e"),
  2265 => (x"4f",x"26",x"48",x"bf"),
  2266 => (x"c4",x"4a",x"71",x"1e"),
  2267 => (x"49",x"72",x"1e",x"66"),
  2268 => (x"26",x"87",x"c1",x"e9"),
  2269 => (x"c2",x"1e",x"4f",x"26"),
  2270 => (x"49",x"bf",x"c3",x"da"),
  2271 => (x"87",x"dc",x"d2",x"c1"),
  2272 => (x"48",x"d2",x"c1",x"c4"),
  2273 => (x"c4",x"78",x"bf",x"e8"),
  2274 => (x"ec",x"48",x"ce",x"c1"),
  2275 => (x"c1",x"c4",x"78",x"bf"),
  2276 => (x"49",x"4a",x"bf",x"d2"),
  2277 => (x"c8",x"99",x"ff",x"c3"),
  2278 => (x"48",x"72",x"2a",x"b7"),
  2279 => (x"c1",x"c4",x"b0",x"71"),
  2280 => (x"4f",x"26",x"58",x"da"),
  2281 => (x"5c",x"5b",x"5e",x"0e"),
  2282 => (x"4b",x"71",x"0e",x"5d"),
  2283 => (x"c4",x"87",x"c7",x"ff"),
  2284 => (x"c0",x"48",x"cd",x"c1"),
  2285 => (x"e5",x"49",x"73",x"50"),
  2286 => (x"49",x"70",x"87",x"c0"),
  2287 => (x"cb",x"9c",x"c2",x"4c"),
  2288 => (x"c6",x"cb",x"49",x"ee"),
  2289 => (x"4d",x"49",x"70",x"87"),
  2290 => (x"97",x"cd",x"c1",x"c4"),
  2291 => (x"e2",x"c1",x"05",x"bf"),
  2292 => (x"49",x"66",x"d0",x"87"),
  2293 => (x"bf",x"d6",x"c1",x"c4"),
  2294 => (x"87",x"d6",x"05",x"99"),
  2295 => (x"c4",x"49",x"66",x"d4"),
  2296 => (x"99",x"bf",x"ce",x"c1"),
  2297 => (x"73",x"87",x"cb",x"05"),
  2298 => (x"87",x"ce",x"e4",x"49"),
  2299 => (x"c1",x"02",x"98",x"70"),
  2300 => (x"4c",x"c1",x"87",x"c1"),
  2301 => (x"75",x"87",x"ff",x"fd"),
  2302 => (x"87",x"db",x"ca",x"49"),
  2303 => (x"c6",x"02",x"98",x"70"),
  2304 => (x"cd",x"c1",x"c4",x"87"),
  2305 => (x"c4",x"50",x"c1",x"48"),
  2306 => (x"bf",x"97",x"cd",x"c1"),
  2307 => (x"87",x"e3",x"c0",x"05"),
  2308 => (x"bf",x"d6",x"c1",x"c4"),
  2309 => (x"99",x"66",x"d0",x"49"),
  2310 => (x"87",x"d6",x"ff",x"05"),
  2311 => (x"bf",x"ce",x"c1",x"c4"),
  2312 => (x"99",x"66",x"d4",x"49"),
  2313 => (x"87",x"ca",x"ff",x"05"),
  2314 => (x"cd",x"e3",x"49",x"73"),
  2315 => (x"05",x"98",x"70",x"87"),
  2316 => (x"74",x"87",x"ff",x"fe"),
  2317 => (x"87",x"d3",x"fb",x"48"),
  2318 => (x"5c",x"5b",x"5e",x"0e"),
  2319 => (x"86",x"f4",x"0e",x"5d"),
  2320 => (x"ec",x"4c",x"4d",x"c0"),
  2321 => (x"a6",x"c4",x"7e",x"bf"),
  2322 => (x"da",x"c1",x"c4",x"48"),
  2323 => (x"1e",x"c1",x"78",x"bf"),
  2324 => (x"d8",x"c1",x"1e",x"c0"),
  2325 => (x"87",x"cc",x"fd",x"49"),
  2326 => (x"98",x"70",x"86",x"c8"),
  2327 => (x"ff",x"87",x"cc",x"02"),
  2328 => (x"87",x"c2",x"fb",x"49"),
  2329 => (x"d1",x"e2",x"49",x"dc"),
  2330 => (x"c4",x"4d",x"c1",x"87"),
  2331 => (x"bf",x"97",x"cd",x"c1"),
  2332 => (x"c0",x"87",x"c4",x"02"),
  2333 => (x"c4",x"87",x"e4",x"fd"),
  2334 => (x"4b",x"bf",x"d2",x"c1"),
  2335 => (x"bf",x"c3",x"da",x"c2"),
  2336 => (x"87",x"e9",x"c0",x"05"),
  2337 => (x"e1",x"49",x"c9",x"c3"),
  2338 => (x"e1",x"c3",x"87",x"f0"),
  2339 => (x"87",x"ea",x"e1",x"49"),
  2340 => (x"ff",x"c3",x"49",x"73"),
  2341 => (x"c0",x"1e",x"71",x"99"),
  2342 => (x"87",x"cc",x"fb",x"49"),
  2343 => (x"b7",x"c8",x"49",x"73"),
  2344 => (x"c1",x"1e",x"71",x"29"),
  2345 => (x"87",x"c0",x"fb",x"49"),
  2346 => (x"fc",x"c5",x"86",x"c8"),
  2347 => (x"d6",x"c1",x"c4",x"87"),
  2348 => (x"02",x"9b",x"4b",x"bf"),
  2349 => (x"d9",x"c2",x"87",x"dd"),
  2350 => (x"c7",x"49",x"bf",x"ff"),
  2351 => (x"98",x"70",x"87",x"d9"),
  2352 => (x"c0",x"87",x"c4",x"05"),
  2353 => (x"c2",x"87",x"d2",x"4b"),
  2354 => (x"fe",x"c6",x"49",x"e0"),
  2355 => (x"c3",x"da",x"c2",x"87"),
  2356 => (x"c2",x"87",x"c6",x"58"),
  2357 => (x"c0",x"48",x"ff",x"d9"),
  2358 => (x"c2",x"49",x"73",x"78"),
  2359 => (x"87",x"cd",x"05",x"99"),
  2360 => (x"e0",x"49",x"cb",x"c3"),
  2361 => (x"49",x"70",x"87",x"d4"),
  2362 => (x"c2",x"02",x"99",x"c2"),
  2363 => (x"73",x"4c",x"fb",x"87"),
  2364 => (x"05",x"99",x"c1",x"49"),
  2365 => (x"cd",x"c3",x"87",x"ce"),
  2366 => (x"fd",x"df",x"ff",x"49"),
  2367 => (x"c2",x"49",x"70",x"87"),
  2368 => (x"87",x"c2",x"02",x"99"),
  2369 => (x"49",x"73",x"4c",x"fa"),
  2370 => (x"ce",x"05",x"99",x"c8"),
  2371 => (x"49",x"c8",x"c3",x"87"),
  2372 => (x"87",x"e6",x"df",x"ff"),
  2373 => (x"99",x"c2",x"49",x"70"),
  2374 => (x"c4",x"87",x"d5",x"02"),
  2375 => (x"02",x"bf",x"de",x"c1"),
  2376 => (x"c1",x"48",x"87",x"ca"),
  2377 => (x"e2",x"c1",x"c4",x"88"),
  2378 => (x"87",x"c2",x"c0",x"58"),
  2379 => (x"4d",x"c1",x"4c",x"ff"),
  2380 => (x"99",x"c4",x"49",x"73"),
  2381 => (x"c3",x"87",x"ce",x"05"),
  2382 => (x"de",x"ff",x"49",x"d0"),
  2383 => (x"49",x"70",x"87",x"fc"),
  2384 => (x"db",x"02",x"99",x"c2"),
  2385 => (x"de",x"c1",x"c4",x"87"),
  2386 => (x"c7",x"48",x"7e",x"bf"),
  2387 => (x"cb",x"03",x"a8",x"b7"),
  2388 => (x"c1",x"48",x"6e",x"87"),
  2389 => (x"e2",x"c1",x"c4",x"80"),
  2390 => (x"87",x"c2",x"c0",x"58"),
  2391 => (x"4d",x"c1",x"4c",x"fe"),
  2392 => (x"ff",x"49",x"c9",x"c3"),
  2393 => (x"70",x"87",x"d3",x"de"),
  2394 => (x"02",x"99",x"c2",x"49"),
  2395 => (x"c1",x"c4",x"87",x"d5"),
  2396 => (x"c0",x"02",x"bf",x"de"),
  2397 => (x"c1",x"c4",x"87",x"c9"),
  2398 => (x"78",x"c0",x"48",x"de"),
  2399 => (x"fd",x"87",x"c2",x"c0"),
  2400 => (x"c3",x"4d",x"c1",x"4c"),
  2401 => (x"dd",x"ff",x"49",x"e1"),
  2402 => (x"49",x"70",x"87",x"f0"),
  2403 => (x"d9",x"02",x"99",x"c2"),
  2404 => (x"de",x"c1",x"c4",x"87"),
  2405 => (x"b7",x"c7",x"48",x"bf"),
  2406 => (x"c9",x"c0",x"03",x"a8"),
  2407 => (x"de",x"c1",x"c4",x"87"),
  2408 => (x"c0",x"78",x"c7",x"48"),
  2409 => (x"4c",x"fc",x"87",x"c2"),
  2410 => (x"b7",x"c0",x"4d",x"c1"),
  2411 => (x"d1",x"c0",x"03",x"ac"),
  2412 => (x"4a",x"66",x"c4",x"87"),
  2413 => (x"6a",x"82",x"d8",x"c1"),
  2414 => (x"87",x"c6",x"c0",x"02"),
  2415 => (x"49",x"74",x"4b",x"6a"),
  2416 => (x"1e",x"c0",x"0f",x"73"),
  2417 => (x"dc",x"1e",x"f0",x"c3"),
  2418 => (x"87",x"d8",x"f7",x"49"),
  2419 => (x"98",x"70",x"86",x"c8"),
  2420 => (x"87",x"e2",x"c0",x"02"),
  2421 => (x"c4",x"48",x"a6",x"c8"),
  2422 => (x"78",x"bf",x"de",x"c1"),
  2423 => (x"cb",x"49",x"66",x"c8"),
  2424 => (x"48",x"66",x"c4",x"91"),
  2425 => (x"7e",x"70",x"80",x"71"),
  2426 => (x"c0",x"02",x"bf",x"6e"),
  2427 => (x"bf",x"6e",x"87",x"c8"),
  2428 => (x"49",x"66",x"c8",x"4b"),
  2429 => (x"9d",x"75",x"0f",x"73"),
  2430 => (x"87",x"c8",x"c0",x"02"),
  2431 => (x"bf",x"de",x"c1",x"c4"),
  2432 => (x"87",x"fd",x"f2",x"49"),
  2433 => (x"bf",x"c7",x"da",x"c2"),
  2434 => (x"87",x"dd",x"c0",x"02"),
  2435 => (x"87",x"c7",x"c2",x"49"),
  2436 => (x"c0",x"02",x"98",x"70"),
  2437 => (x"c1",x"c4",x"87",x"d3"),
  2438 => (x"f2",x"49",x"bf",x"de"),
  2439 => (x"49",x"c0",x"87",x"e3"),
  2440 => (x"c2",x"87",x"c3",x"f4"),
  2441 => (x"c0",x"48",x"c7",x"da"),
  2442 => (x"f3",x"8e",x"f4",x"78"),
  2443 => (x"5e",x"0e",x"87",x"dd"),
  2444 => (x"0e",x"5d",x"5c",x"5b"),
  2445 => (x"c4",x"4c",x"71",x"1e"),
  2446 => (x"49",x"bf",x"da",x"c1"),
  2447 => (x"4d",x"a1",x"cd",x"c1"),
  2448 => (x"69",x"81",x"d1",x"c1"),
  2449 => (x"02",x"9c",x"74",x"7e"),
  2450 => (x"a5",x"c4",x"87",x"cf"),
  2451 => (x"c4",x"7b",x"74",x"4b"),
  2452 => (x"49",x"bf",x"da",x"c1"),
  2453 => (x"6e",x"87",x"fc",x"f2"),
  2454 => (x"05",x"9c",x"74",x"7b"),
  2455 => (x"4b",x"c0",x"87",x"c4"),
  2456 => (x"4b",x"c1",x"87",x"c2"),
  2457 => (x"fd",x"f2",x"49",x"73"),
  2458 => (x"02",x"66",x"d4",x"87"),
  2459 => (x"da",x"49",x"87",x"c7"),
  2460 => (x"c2",x"4a",x"70",x"87"),
  2461 => (x"c2",x"4a",x"c0",x"87"),
  2462 => (x"26",x"5a",x"cb",x"da"),
  2463 => (x"00",x"87",x"cc",x"f2"),
  2464 => (x"00",x"00",x"00",x"00"),
  2465 => (x"00",x"00",x"00",x"00"),
  2466 => (x"1e",x"00",x"00",x"00"),
  2467 => (x"c8",x"ff",x"4a",x"71"),
  2468 => (x"a1",x"72",x"49",x"bf"),
  2469 => (x"1e",x"4f",x"26",x"48"),
  2470 => (x"89",x"bf",x"c8",x"ff"),
  2471 => (x"c0",x"c0",x"c0",x"fe"),
  2472 => (x"01",x"a9",x"c0",x"c0"),
  2473 => (x"4a",x"c0",x"87",x"c4"),
  2474 => (x"4a",x"c1",x"87",x"c2"),
  2475 => (x"4f",x"26",x"48",x"72"),
  2476 => (x"5c",x"5b",x"5e",x"0e"),
  2477 => (x"4b",x"71",x"0e",x"5d"),
  2478 => (x"d0",x"4c",x"d4",x"ff"),
  2479 => (x"78",x"c0",x"48",x"66"),
  2480 => (x"da",x"ff",x"49",x"d6"),
  2481 => (x"ff",x"c3",x"87",x"f4"),
  2482 => (x"c3",x"49",x"6c",x"7c"),
  2483 => (x"4d",x"71",x"99",x"ff"),
  2484 => (x"99",x"f0",x"c3",x"49"),
  2485 => (x"05",x"a9",x"e0",x"c1"),
  2486 => (x"ff",x"c3",x"87",x"cb"),
  2487 => (x"c3",x"48",x"6c",x"7c"),
  2488 => (x"08",x"66",x"d0",x"98"),
  2489 => (x"7c",x"ff",x"c3",x"78"),
  2490 => (x"c8",x"49",x"4a",x"6c"),
  2491 => (x"7c",x"ff",x"c3",x"31"),
  2492 => (x"b2",x"71",x"4a",x"6c"),
  2493 => (x"31",x"c8",x"49",x"72"),
  2494 => (x"6c",x"7c",x"ff",x"c3"),
  2495 => (x"72",x"b2",x"71",x"4a"),
  2496 => (x"c3",x"31",x"c8",x"49"),
  2497 => (x"4a",x"6c",x"7c",x"ff"),
  2498 => (x"d0",x"ff",x"b2",x"71"),
  2499 => (x"78",x"e0",x"c0",x"48"),
  2500 => (x"c2",x"02",x"9b",x"73"),
  2501 => (x"75",x"7b",x"72",x"87"),
  2502 => (x"26",x"4d",x"26",x"48"),
  2503 => (x"26",x"4b",x"26",x"4c"),
  2504 => (x"4f",x"26",x"1e",x"4f"),
  2505 => (x"5c",x"5b",x"5e",x"0e"),
  2506 => (x"76",x"86",x"f8",x"0e"),
  2507 => (x"49",x"a6",x"c8",x"1e"),
  2508 => (x"c4",x"87",x"fd",x"fd"),
  2509 => (x"6e",x"4b",x"70",x"86"),
  2510 => (x"03",x"a8",x"c2",x"48"),
  2511 => (x"73",x"87",x"ca",x"c3"),
  2512 => (x"9a",x"f0",x"c3",x"4a"),
  2513 => (x"02",x"aa",x"d0",x"c1"),
  2514 => (x"e0",x"c1",x"87",x"c7"),
  2515 => (x"f8",x"c2",x"05",x"aa"),
  2516 => (x"c8",x"49",x"73",x"87"),
  2517 => (x"87",x"c3",x"02",x"99"),
  2518 => (x"73",x"87",x"c6",x"ff"),
  2519 => (x"c2",x"9c",x"c3",x"4c"),
  2520 => (x"cf",x"c1",x"05",x"ac"),
  2521 => (x"49",x"66",x"c4",x"87"),
  2522 => (x"1e",x"71",x"31",x"c9"),
  2523 => (x"c2",x"4a",x"66",x"c4"),
  2524 => (x"c1",x"c4",x"92",x"d8"),
  2525 => (x"81",x"72",x"49",x"e2"),
  2526 => (x"87",x"c2",x"d0",x"fe"),
  2527 => (x"1e",x"49",x"66",x"c4"),
  2528 => (x"ff",x"49",x"e3",x"c0"),
  2529 => (x"d8",x"87",x"d8",x"d8"),
  2530 => (x"ed",x"d7",x"ff",x"49"),
  2531 => (x"1e",x"c0",x"c8",x"87"),
  2532 => (x"49",x"d2",x"f0",x"c3"),
  2533 => (x"87",x"f3",x"e7",x"fd"),
  2534 => (x"c0",x"48",x"d0",x"ff"),
  2535 => (x"f0",x"c3",x"78",x"e0"),
  2536 => (x"66",x"d0",x"1e",x"d2"),
  2537 => (x"92",x"d8",x"c2",x"4a"),
  2538 => (x"49",x"e2",x"c1",x"c4"),
  2539 => (x"ca",x"fe",x"81",x"72"),
  2540 => (x"86",x"d0",x"87",x"dd"),
  2541 => (x"c1",x"05",x"ac",x"c1"),
  2542 => (x"66",x"c4",x"87",x"cf"),
  2543 => (x"71",x"31",x"c9",x"49"),
  2544 => (x"4a",x"66",x"c4",x"1e"),
  2545 => (x"c4",x"92",x"d8",x"c2"),
  2546 => (x"72",x"49",x"e2",x"c1"),
  2547 => (x"ed",x"ce",x"fe",x"81"),
  2548 => (x"d2",x"f0",x"c3",x"87"),
  2549 => (x"4a",x"66",x"c8",x"1e"),
  2550 => (x"c4",x"92",x"d8",x"c2"),
  2551 => (x"72",x"49",x"e2",x"c1"),
  2552 => (x"e7",x"c8",x"fe",x"81"),
  2553 => (x"49",x"66",x"c8",x"87"),
  2554 => (x"49",x"e3",x"c0",x"1e"),
  2555 => (x"87",x"ef",x"d6",x"ff"),
  2556 => (x"d6",x"ff",x"49",x"d7"),
  2557 => (x"c0",x"c8",x"87",x"c4"),
  2558 => (x"d2",x"f0",x"c3",x"1e"),
  2559 => (x"f4",x"e5",x"fd",x"49"),
  2560 => (x"ff",x"86",x"d0",x"87"),
  2561 => (x"e0",x"c0",x"48",x"d0"),
  2562 => (x"fc",x"8e",x"f8",x"78"),
  2563 => (x"5e",x"0e",x"87",x"cd"),
  2564 => (x"0e",x"5d",x"5c",x"5b"),
  2565 => (x"ff",x"4d",x"71",x"1e"),
  2566 => (x"66",x"d4",x"4c",x"d4"),
  2567 => (x"b7",x"c3",x"48",x"7e"),
  2568 => (x"87",x"c5",x"06",x"a8"),
  2569 => (x"e3",x"c1",x"48",x"c0"),
  2570 => (x"fe",x"49",x"75",x"87"),
  2571 => (x"75",x"87",x"f7",x"df"),
  2572 => (x"4b",x"66",x"c4",x"1e"),
  2573 => (x"c4",x"93",x"d8",x"c2"),
  2574 => (x"73",x"83",x"e2",x"c1"),
  2575 => (x"fe",x"c2",x"fe",x"49"),
  2576 => (x"6b",x"83",x"c8",x"87"),
  2577 => (x"48",x"d0",x"ff",x"4b"),
  2578 => (x"dd",x"78",x"e1",x"c8"),
  2579 => (x"c3",x"49",x"73",x"7c"),
  2580 => (x"7c",x"71",x"99",x"ff"),
  2581 => (x"b7",x"c8",x"49",x"73"),
  2582 => (x"99",x"ff",x"c3",x"29"),
  2583 => (x"49",x"73",x"7c",x"71"),
  2584 => (x"c3",x"29",x"b7",x"d0"),
  2585 => (x"7c",x"71",x"99",x"ff"),
  2586 => (x"b7",x"d8",x"49",x"73"),
  2587 => (x"c0",x"7c",x"71",x"29"),
  2588 => (x"7c",x"7c",x"7c",x"7c"),
  2589 => (x"7c",x"7c",x"7c",x"7c"),
  2590 => (x"7c",x"7c",x"7c",x"7c"),
  2591 => (x"c4",x"78",x"e0",x"c0"),
  2592 => (x"49",x"dc",x"1e",x"66"),
  2593 => (x"87",x"d7",x"d4",x"ff"),
  2594 => (x"48",x"73",x"86",x"c8"),
  2595 => (x"87",x"c9",x"fa",x"26"),
  2596 => (x"4a",x"d4",x"ff",x"1e"),
  2597 => (x"c8",x"48",x"d0",x"ff"),
  2598 => (x"f0",x"c3",x"78",x"c5"),
  2599 => (x"c0",x"7a",x"71",x"7a"),
  2600 => (x"7a",x"7a",x"7a",x"7a"),
  2601 => (x"4f",x"26",x"78",x"c4"),
  2602 => (x"4a",x"d4",x"ff",x"1e"),
  2603 => (x"c8",x"48",x"d0",x"ff"),
  2604 => (x"7a",x"c0",x"78",x"c5"),
  2605 => (x"7a",x"c0",x"49",x"6a"),
  2606 => (x"7a",x"7a",x"7a",x"7a"),
  2607 => (x"48",x"71",x"78",x"c4"),
  2608 => (x"5e",x"0e",x"4f",x"26"),
  2609 => (x"0e",x"5d",x"5c",x"5b"),
  2610 => (x"a6",x"cc",x"86",x"e4"),
  2611 => (x"66",x"ec",x"c0",x"59"),
  2612 => (x"58",x"a6",x"dc",x"48"),
  2613 => (x"e8",x"c2",x"4d",x"70"),
  2614 => (x"d2",x"c6",x"c4",x"95"),
  2615 => (x"a5",x"d8",x"c2",x"85"),
  2616 => (x"48",x"a6",x"c4",x"7e"),
  2617 => (x"78",x"a5",x"dc",x"c2"),
  2618 => (x"4c",x"bf",x"66",x"c4"),
  2619 => (x"c2",x"94",x"bf",x"6e"),
  2620 => (x"94",x"6d",x"85",x"e0"),
  2621 => (x"c0",x"4b",x"66",x"c8"),
  2622 => (x"49",x"c0",x"c8",x"4a"),
  2623 => (x"87",x"c3",x"e0",x"fd"),
  2624 => (x"c1",x"48",x"66",x"c8"),
  2625 => (x"c8",x"78",x"9f",x"c0"),
  2626 => (x"81",x"c2",x"49",x"66"),
  2627 => (x"79",x"9f",x"bf",x"6e"),
  2628 => (x"c6",x"49",x"66",x"c8"),
  2629 => (x"bf",x"66",x"c4",x"81"),
  2630 => (x"66",x"c8",x"79",x"9f"),
  2631 => (x"6d",x"81",x"cc",x"49"),
  2632 => (x"66",x"c8",x"79",x"9f"),
  2633 => (x"d0",x"80",x"d4",x"48"),
  2634 => (x"e7",x"c2",x"58",x"a6"),
  2635 => (x"66",x"cc",x"48",x"fb"),
  2636 => (x"4a",x"a1",x"d4",x"49"),
  2637 => (x"aa",x"71",x"41",x"20"),
  2638 => (x"c8",x"87",x"f9",x"05"),
  2639 => (x"ee",x"c0",x"48",x"66"),
  2640 => (x"58",x"a6",x"d4",x"80"),
  2641 => (x"48",x"d0",x"e8",x"c2"),
  2642 => (x"c8",x"49",x"66",x"d0"),
  2643 => (x"41",x"20",x"4a",x"a1"),
  2644 => (x"f9",x"05",x"aa",x"71"),
  2645 => (x"48",x"66",x"c8",x"87"),
  2646 => (x"d8",x"80",x"f6",x"c0"),
  2647 => (x"e8",x"c2",x"58",x"a6"),
  2648 => (x"66",x"d4",x"48",x"d9"),
  2649 => (x"a1",x"e8",x"c0",x"49"),
  2650 => (x"71",x"41",x"20",x"4a"),
  2651 => (x"87",x"f9",x"05",x"aa"),
  2652 => (x"c0",x"4a",x"66",x"d8"),
  2653 => (x"66",x"d4",x"82",x"f1"),
  2654 => (x"72",x"81",x"cb",x"49"),
  2655 => (x"49",x"66",x"c8",x"51"),
  2656 => (x"c8",x"81",x"de",x"c1"),
  2657 => (x"79",x"9f",x"d0",x"c0"),
  2658 => (x"c1",x"49",x"66",x"c8"),
  2659 => (x"c0",x"c8",x"81",x"e2"),
  2660 => (x"66",x"c8",x"79",x"9f"),
  2661 => (x"81",x"ea",x"c1",x"49"),
  2662 => (x"c8",x"79",x"9f",x"c1"),
  2663 => (x"ec",x"c1",x"49",x"66"),
  2664 => (x"9f",x"bf",x"6e",x"81"),
  2665 => (x"49",x"66",x"c8",x"79"),
  2666 => (x"c4",x"81",x"ee",x"c1"),
  2667 => (x"79",x"9f",x"bf",x"66"),
  2668 => (x"c1",x"49",x"66",x"c8"),
  2669 => (x"9f",x"6d",x"81",x"f0"),
  2670 => (x"cf",x"4b",x"74",x"79"),
  2671 => (x"73",x"9b",x"ff",x"ff"),
  2672 => (x"49",x"66",x"c8",x"4a"),
  2673 => (x"72",x"81",x"f2",x"c1"),
  2674 => (x"4a",x"74",x"79",x"9f"),
  2675 => (x"ff",x"cf",x"2a",x"d0"),
  2676 => (x"4c",x"72",x"9a",x"ff"),
  2677 => (x"c1",x"49",x"66",x"c8"),
  2678 => (x"9f",x"74",x"81",x"f4"),
  2679 => (x"66",x"c8",x"73",x"79"),
  2680 => (x"81",x"f8",x"c1",x"49"),
  2681 => (x"72",x"79",x"9f",x"73"),
  2682 => (x"c1",x"49",x"66",x"c8"),
  2683 => (x"9f",x"72",x"81",x"fa"),
  2684 => (x"26",x"8e",x"e4",x"79"),
  2685 => (x"26",x"4c",x"26",x"4d"),
  2686 => (x"69",x"4f",x"26",x"4b"),
  2687 => (x"69",x"53",x"54",x"4d"),
  2688 => (x"69",x"6e",x"69",x"4d"),
  2689 => (x"72",x"67",x"48",x"4d"),
  2690 => (x"6c",x"64",x"66",x"61"),
  2691 => (x"00",x"65",x"20",x"69"),
  2692 => (x"30",x"30",x"31",x"2e"),
  2693 => (x"20",x"20",x"20",x"20"),
  2694 => (x"69",x"44",x"65",x"00"),
  2695 => (x"66",x"53",x"54",x"4d"),
  2696 => (x"20",x"79",x"20",x"69"),
  2697 => (x"20",x"20",x"20",x"20"),
  2698 => (x"20",x"20",x"20",x"20"),
  2699 => (x"20",x"20",x"20",x"20"),
  2700 => (x"20",x"20",x"20",x"20"),
  2701 => (x"20",x"20",x"20",x"20"),
  2702 => (x"20",x"20",x"20",x"20"),
  2703 => (x"20",x"20",x"20",x"20"),
  2704 => (x"73",x"1e",x"00",x"20"),
  2705 => (x"d4",x"4b",x"71",x"1e"),
  2706 => (x"87",x"d4",x"02",x"66"),
  2707 => (x"d8",x"49",x"66",x"c8"),
  2708 => (x"c8",x"4a",x"73",x"31"),
  2709 => (x"49",x"a1",x"72",x"32"),
  2710 => (x"71",x"81",x"66",x"cc"),
  2711 => (x"87",x"e3",x"c0",x"48"),
  2712 => (x"c2",x"49",x"66",x"d0"),
  2713 => (x"c6",x"c4",x"91",x"e8"),
  2714 => (x"dc",x"c2",x"81",x"d2"),
  2715 => (x"4a",x"6a",x"4a",x"a1"),
  2716 => (x"66",x"c8",x"92",x"73"),
  2717 => (x"81",x"e0",x"c2",x"82"),
  2718 => (x"91",x"72",x"49",x"69"),
  2719 => (x"c1",x"81",x"66",x"cc"),
  2720 => (x"fd",x"48",x"71",x"89"),
  2721 => (x"71",x"1e",x"87",x"f1"),
  2722 => (x"49",x"d4",x"ff",x"4a"),
  2723 => (x"c8",x"48",x"d0",x"ff"),
  2724 => (x"d0",x"c2",x"78",x"c5"),
  2725 => (x"79",x"79",x"c0",x"79"),
  2726 => (x"79",x"79",x"79",x"79"),
  2727 => (x"79",x"72",x"79",x"79"),
  2728 => (x"66",x"c4",x"79",x"c0"),
  2729 => (x"c8",x"79",x"c0",x"79"),
  2730 => (x"79",x"c0",x"79",x"66"),
  2731 => (x"c0",x"79",x"66",x"cc"),
  2732 => (x"79",x"66",x"d0",x"79"),
  2733 => (x"66",x"d4",x"79",x"c0"),
  2734 => (x"26",x"78",x"c4",x"79"),
  2735 => (x"4a",x"71",x"1e",x"4f"),
  2736 => (x"97",x"49",x"a2",x"c6"),
  2737 => (x"f0",x"c3",x"49",x"69"),
  2738 => (x"c0",x"1e",x"71",x"99"),
  2739 => (x"1e",x"c1",x"1e",x"1e"),
  2740 => (x"fe",x"49",x"1e",x"c0"),
  2741 => (x"d0",x"c2",x"87",x"f0"),
  2742 => (x"87",x"f4",x"f6",x"49"),
  2743 => (x"4f",x"26",x"8e",x"ec"),
  2744 => (x"1e",x"1e",x"c0",x"1e"),
  2745 => (x"c1",x"1e",x"1e",x"1e"),
  2746 => (x"87",x"da",x"fe",x"49"),
  2747 => (x"f6",x"49",x"d0",x"c2"),
  2748 => (x"8e",x"ec",x"87",x"de"),
  2749 => (x"71",x"1e",x"4f",x"26"),
  2750 => (x"48",x"d0",x"ff",x"4a"),
  2751 => (x"ff",x"78",x"c5",x"c8"),
  2752 => (x"e0",x"c2",x"48",x"d4"),
  2753 => (x"78",x"78",x"c0",x"78"),
  2754 => (x"c8",x"78",x"78",x"78"),
  2755 => (x"49",x"72",x"1e",x"c0"),
  2756 => (x"87",x"e1",x"d9",x"fd"),
  2757 => (x"c4",x"48",x"d0",x"ff"),
  2758 => (x"4f",x"26",x"26",x"78"),
  2759 => (x"5c",x"5b",x"5e",x"0e"),
  2760 => (x"86",x"f8",x"0e",x"5d"),
  2761 => (x"a2",x"c2",x"4a",x"71"),
  2762 => (x"7b",x"97",x"c1",x"4b"),
  2763 => (x"c1",x"4c",x"a2",x"c3"),
  2764 => (x"49",x"a2",x"7c",x"97"),
  2765 => (x"a2",x"c4",x"51",x"c0"),
  2766 => (x"7d",x"97",x"c0",x"4d"),
  2767 => (x"6e",x"7e",x"a2",x"c5"),
  2768 => (x"c4",x"50",x"c0",x"48"),
  2769 => (x"a2",x"c6",x"48",x"a6"),
  2770 => (x"48",x"66",x"c4",x"78"),
  2771 => (x"66",x"d8",x"50",x"c0"),
  2772 => (x"d2",x"f0",x"c3",x"1e"),
  2773 => (x"87",x"ea",x"f5",x"49"),
  2774 => (x"bf",x"97",x"66",x"c8"),
  2775 => (x"66",x"c8",x"1e",x"49"),
  2776 => (x"1e",x"49",x"bf",x"97"),
  2777 => (x"14",x"1e",x"49",x"15"),
  2778 => (x"49",x"13",x"1e",x"49"),
  2779 => (x"fc",x"49",x"c0",x"1e"),
  2780 => (x"49",x"c8",x"87",x"d4"),
  2781 => (x"c3",x"87",x"d9",x"f4"),
  2782 => (x"fd",x"49",x"d2",x"f0"),
  2783 => (x"49",x"d0",x"87",x"f8"),
  2784 => (x"e0",x"87",x"cd",x"f4"),
  2785 => (x"87",x"eb",x"f9",x"8e"),
  2786 => (x"c6",x"4a",x"71",x"1e"),
  2787 => (x"69",x"97",x"49",x"a2"),
  2788 => (x"a2",x"c5",x"1e",x"49"),
  2789 => (x"49",x"69",x"97",x"49"),
  2790 => (x"49",x"a2",x"c4",x"1e"),
  2791 => (x"1e",x"49",x"69",x"97"),
  2792 => (x"97",x"49",x"a2",x"c3"),
  2793 => (x"c2",x"1e",x"49",x"69"),
  2794 => (x"69",x"97",x"49",x"a2"),
  2795 => (x"49",x"c0",x"1e",x"49"),
  2796 => (x"c2",x"87",x"d3",x"fb"),
  2797 => (x"d7",x"f3",x"49",x"d0"),
  2798 => (x"26",x"8e",x"ec",x"87"),
  2799 => (x"1e",x"73",x"1e",x"4f"),
  2800 => (x"a2",x"c2",x"4a",x"71"),
  2801 => (x"d0",x"4b",x"11",x"49"),
  2802 => (x"c8",x"06",x"ab",x"b7"),
  2803 => (x"49",x"d1",x"c2",x"87"),
  2804 => (x"d5",x"87",x"fd",x"f2"),
  2805 => (x"49",x"66",x"c8",x"87"),
  2806 => (x"c4",x"91",x"e8",x"c2"),
  2807 => (x"c2",x"81",x"d2",x"c6"),
  2808 => (x"79",x"73",x"81",x"e4"),
  2809 => (x"f2",x"49",x"d0",x"c2"),
  2810 => (x"ca",x"f8",x"87",x"e6"),
  2811 => (x"1e",x"73",x"1e",x"87"),
  2812 => (x"a3",x"c6",x"4b",x"71"),
  2813 => (x"49",x"69",x"97",x"49"),
  2814 => (x"49",x"a3",x"c5",x"1e"),
  2815 => (x"1e",x"49",x"69",x"97"),
  2816 => (x"97",x"49",x"a3",x"c4"),
  2817 => (x"c3",x"1e",x"49",x"69"),
  2818 => (x"69",x"97",x"49",x"a3"),
  2819 => (x"a3",x"c2",x"1e",x"49"),
  2820 => (x"49",x"69",x"97",x"49"),
  2821 => (x"4a",x"a3",x"c1",x"1e"),
  2822 => (x"e9",x"f9",x"49",x"12"),
  2823 => (x"49",x"d0",x"c2",x"87"),
  2824 => (x"ec",x"87",x"ed",x"f1"),
  2825 => (x"87",x"cf",x"f7",x"8e"),
  2826 => (x"5c",x"5b",x"5e",x"0e"),
  2827 => (x"71",x"1e",x"0e",x"5d"),
  2828 => (x"c2",x"49",x"6e",x"7e"),
  2829 => (x"79",x"97",x"c1",x"81"),
  2830 => (x"83",x"c3",x"4b",x"6e"),
  2831 => (x"6e",x"7b",x"97",x"c1"),
  2832 => (x"c0",x"82",x"c1",x"4a"),
  2833 => (x"4c",x"6e",x"7a",x"97"),
  2834 => (x"97",x"c0",x"84",x"c4"),
  2835 => (x"c5",x"4d",x"6e",x"7c"),
  2836 => (x"6e",x"55",x"c0",x"85"),
  2837 => (x"97",x"85",x"c6",x"4d"),
  2838 => (x"c0",x"1e",x"4d",x"6d"),
  2839 => (x"4c",x"6c",x"97",x"1e"),
  2840 => (x"4b",x"6b",x"97",x"1e"),
  2841 => (x"49",x"69",x"97",x"1e"),
  2842 => (x"f8",x"49",x"12",x"1e"),
  2843 => (x"d0",x"c2",x"87",x"d8"),
  2844 => (x"87",x"dc",x"f0",x"49"),
  2845 => (x"fa",x"f5",x"8e",x"e8"),
  2846 => (x"5b",x"5e",x"0e",x"87"),
  2847 => (x"ff",x"0e",x"5d",x"5c"),
  2848 => (x"4c",x"71",x"86",x"dc"),
  2849 => (x"11",x"49",x"a4",x"c3"),
  2850 => (x"4a",x"a4",x"c4",x"4d"),
  2851 => (x"97",x"49",x"a4",x"c5"),
  2852 => (x"31",x"c8",x"49",x"69"),
  2853 => (x"48",x"4a",x"6a",x"97"),
  2854 => (x"a6",x"d4",x"b0",x"71"),
  2855 => (x"7e",x"a4",x"c6",x"58"),
  2856 => (x"49",x"bf",x"97",x"6e"),
  2857 => (x"d8",x"98",x"cf",x"48"),
  2858 => (x"48",x"71",x"58",x"a6"),
  2859 => (x"dc",x"98",x"c0",x"c1"),
  2860 => (x"ec",x"48",x"58",x"a6"),
  2861 => (x"78",x"a4",x"c2",x"80"),
  2862 => (x"bf",x"97",x"66",x"c4"),
  2863 => (x"c3",x"05",x"9b",x"4b"),
  2864 => (x"4b",x"c0",x"c4",x"87"),
  2865 => (x"c0",x"1e",x"66",x"d8"),
  2866 => (x"75",x"1e",x"66",x"f8"),
  2867 => (x"66",x"e0",x"c0",x"1e"),
  2868 => (x"66",x"e0",x"c0",x"1e"),
  2869 => (x"87",x"ea",x"f5",x"49"),
  2870 => (x"49",x"70",x"86",x"d0"),
  2871 => (x"59",x"a6",x"e0",x"c0"),
  2872 => (x"c5",x"02",x"9b",x"73"),
  2873 => (x"f8",x"c0",x"87",x"fb"),
  2874 => (x"87",x"c5",x"02",x"66"),
  2875 => (x"c5",x"5b",x"a6",x"d0"),
  2876 => (x"48",x"a6",x"cc",x"87"),
  2877 => (x"66",x"cc",x"78",x"c1"),
  2878 => (x"66",x"f8",x"c0",x"4c"),
  2879 => (x"c0",x"87",x"de",x"02"),
  2880 => (x"c2",x"49",x"66",x"f4"),
  2881 => (x"c6",x"c4",x"91",x"e8"),
  2882 => (x"e4",x"c2",x"81",x"d2"),
  2883 => (x"48",x"a6",x"c8",x"81"),
  2884 => (x"66",x"cc",x"78",x"69"),
  2885 => (x"b7",x"66",x"c8",x"48"),
  2886 => (x"87",x"c1",x"06",x"a8"),
  2887 => (x"66",x"fc",x"c0",x"4c"),
  2888 => (x"c8",x"87",x"d9",x"05"),
  2889 => (x"87",x"e8",x"ed",x"49"),
  2890 => (x"70",x"87",x"fd",x"ed"),
  2891 => (x"05",x"99",x"c4",x"49"),
  2892 => (x"f3",x"ed",x"87",x"ca"),
  2893 => (x"c4",x"49",x"70",x"87"),
  2894 => (x"87",x"f6",x"02",x"99"),
  2895 => (x"88",x"c1",x"48",x"74"),
  2896 => (x"70",x"58",x"a6",x"d0"),
  2897 => (x"02",x"9c",x"74",x"4a"),
  2898 => (x"c1",x"87",x"d4",x"c1"),
  2899 => (x"c2",x"c1",x"02",x"ab"),
  2900 => (x"66",x"f4",x"c0",x"87"),
  2901 => (x"91",x"e8",x"c2",x"49"),
  2902 => (x"48",x"d2",x"c6",x"c4"),
  2903 => (x"a6",x"cc",x"80",x"71"),
  2904 => (x"49",x"66",x"c8",x"58"),
  2905 => (x"69",x"81",x"e0",x"c2"),
  2906 => (x"e4",x"c0",x"05",x"ad"),
  2907 => (x"d4",x"4d",x"c1",x"87"),
  2908 => (x"80",x"c1",x"48",x"66"),
  2909 => (x"c8",x"58",x"a6",x"d8"),
  2910 => (x"dc",x"c2",x"49",x"66"),
  2911 => (x"05",x"a8",x"69",x"81"),
  2912 => (x"a6",x"d4",x"87",x"d1"),
  2913 => (x"d0",x"78",x"c0",x"48"),
  2914 => (x"80",x"c1",x"48",x"66"),
  2915 => (x"c2",x"58",x"a6",x"d4"),
  2916 => (x"c1",x"85",x"c1",x"87"),
  2917 => (x"c1",x"49",x"72",x"8b"),
  2918 => (x"05",x"99",x"71",x"8a"),
  2919 => (x"d8",x"87",x"ec",x"fe"),
  2920 => (x"87",x"d9",x"02",x"66"),
  2921 => (x"66",x"dc",x"49",x"74"),
  2922 => (x"c3",x"4a",x"71",x"81"),
  2923 => (x"4d",x"72",x"9a",x"ff"),
  2924 => (x"b7",x"c8",x"4a",x"71"),
  2925 => (x"5a",x"a6",x"d4",x"2a"),
  2926 => (x"a6",x"29",x"b7",x"d8"),
  2927 => (x"bf",x"97",x"6e",x"59"),
  2928 => (x"99",x"f0",x"c3",x"49"),
  2929 => (x"71",x"b1",x"66",x"d4"),
  2930 => (x"49",x"66",x"d4",x"1e"),
  2931 => (x"71",x"29",x"b7",x"c8"),
  2932 => (x"1e",x"66",x"d8",x"1e"),
  2933 => (x"66",x"d4",x"1e",x"75"),
  2934 => (x"1e",x"49",x"bf",x"97"),
  2935 => (x"e5",x"f2",x"49",x"c0"),
  2936 => (x"c0",x"86",x"d4",x"87"),
  2937 => (x"c1",x"05",x"66",x"fc"),
  2938 => (x"49",x"d0",x"87",x"f1"),
  2939 => (x"c0",x"87",x"e1",x"ea"),
  2940 => (x"c2",x"49",x"66",x"f4"),
  2941 => (x"c6",x"c4",x"91",x"e8"),
  2942 => (x"80",x"71",x"48",x"d2"),
  2943 => (x"c8",x"58",x"a6",x"cc"),
  2944 => (x"81",x"c8",x"49",x"66"),
  2945 => (x"cd",x"c1",x"02",x"69"),
  2946 => (x"49",x"66",x"dc",x"87"),
  2947 => (x"1e",x"71",x"31",x"c9"),
  2948 => (x"fd",x"49",x"66",x"cc"),
  2949 => (x"c4",x"87",x"e7",x"f5"),
  2950 => (x"a6",x"e0",x"c0",x"86"),
  2951 => (x"78",x"66",x"cc",x"48"),
  2952 => (x"c0",x"02",x"9c",x"74"),
  2953 => (x"1e",x"c0",x"87",x"f5"),
  2954 => (x"fd",x"49",x"66",x"cc"),
  2955 => (x"c1",x"87",x"dd",x"ef"),
  2956 => (x"49",x"66",x"d0",x"1e"),
  2957 => (x"87",x"f3",x"ed",x"fd"),
  2958 => (x"66",x"dc",x"86",x"c8"),
  2959 => (x"c0",x"80",x"c1",x"48"),
  2960 => (x"c0",x"58",x"a6",x"e0"),
  2961 => (x"48",x"49",x"66",x"e0"),
  2962 => (x"e4",x"c0",x"88",x"c1"),
  2963 => (x"99",x"71",x"58",x"a6"),
  2964 => (x"87",x"d2",x"ff",x"05"),
  2965 => (x"49",x"c9",x"87",x"c5"),
  2966 => (x"73",x"87",x"f5",x"e8"),
  2967 => (x"c5",x"fa",x"05",x"9b"),
  2968 => (x"66",x"fc",x"c0",x"87"),
  2969 => (x"d0",x"87",x"c5",x"02"),
  2970 => (x"87",x"e4",x"e8",x"49"),
  2971 => (x"ee",x"8e",x"dc",x"ff"),
  2972 => (x"5e",x"0e",x"87",x"c1"),
  2973 => (x"0e",x"5d",x"5c",x"5b"),
  2974 => (x"4c",x"71",x"86",x"e0"),
  2975 => (x"11",x"49",x"a4",x"c3"),
  2976 => (x"58",x"a6",x"d4",x"48"),
  2977 => (x"c5",x"4a",x"a4",x"c4"),
  2978 => (x"69",x"97",x"49",x"a4"),
  2979 => (x"97",x"31",x"c8",x"49"),
  2980 => (x"71",x"48",x"4a",x"6a"),
  2981 => (x"58",x"a6",x"d8",x"b0"),
  2982 => (x"6e",x"7e",x"a4",x"c6"),
  2983 => (x"4d",x"49",x"bf",x"97"),
  2984 => (x"48",x"71",x"9d",x"cf"),
  2985 => (x"dc",x"98",x"c0",x"c1"),
  2986 => (x"ec",x"48",x"58",x"a6"),
  2987 => (x"78",x"a4",x"c2",x"80"),
  2988 => (x"bf",x"97",x"66",x"c4"),
  2989 => (x"1e",x"66",x"d8",x"4b"),
  2990 => (x"1e",x"66",x"f4",x"c0"),
  2991 => (x"75",x"1e",x"66",x"d8"),
  2992 => (x"66",x"e4",x"c0",x"1e"),
  2993 => (x"87",x"fa",x"ed",x"49"),
  2994 => (x"49",x"70",x"86",x"d0"),
  2995 => (x"59",x"a6",x"e0",x"c0"),
  2996 => (x"c3",x"05",x"9b",x"73"),
  2997 => (x"4b",x"c0",x"c4",x"87"),
  2998 => (x"f3",x"e6",x"49",x"c4"),
  2999 => (x"49",x"66",x"dc",x"87"),
  3000 => (x"1e",x"71",x"31",x"c9"),
  3001 => (x"49",x"66",x"f4",x"c0"),
  3002 => (x"c4",x"91",x"e8",x"c2"),
  3003 => (x"71",x"48",x"d2",x"c6"),
  3004 => (x"58",x"a6",x"d4",x"80"),
  3005 => (x"fd",x"49",x"66",x"d0"),
  3006 => (x"c4",x"87",x"c3",x"f2"),
  3007 => (x"02",x"9b",x"73",x"86"),
  3008 => (x"c0",x"87",x"df",x"c4"),
  3009 => (x"c4",x"02",x"66",x"f4"),
  3010 => (x"c2",x"4a",x"73",x"87"),
  3011 => (x"72",x"4a",x"c1",x"87"),
  3012 => (x"66",x"f4",x"c0",x"4c"),
  3013 => (x"cc",x"87",x"d3",x"02"),
  3014 => (x"e4",x"c2",x"49",x"66"),
  3015 => (x"48",x"a6",x"c8",x"81"),
  3016 => (x"66",x"c8",x"78",x"69"),
  3017 => (x"c1",x"06",x"aa",x"b7"),
  3018 => (x"9c",x"74",x"4c",x"87"),
  3019 => (x"87",x"d5",x"c2",x"02"),
  3020 => (x"70",x"87",x"f5",x"e5"),
  3021 => (x"05",x"99",x"c8",x"49"),
  3022 => (x"eb",x"e5",x"87",x"ca"),
  3023 => (x"c8",x"49",x"70",x"87"),
  3024 => (x"87",x"f6",x"02",x"99"),
  3025 => (x"c8",x"48",x"d0",x"ff"),
  3026 => (x"d4",x"ff",x"78",x"c5"),
  3027 => (x"78",x"f0",x"c2",x"48"),
  3028 => (x"78",x"78",x"78",x"c0"),
  3029 => (x"c0",x"c8",x"78",x"78"),
  3030 => (x"d2",x"f0",x"c3",x"1e"),
  3031 => (x"ea",x"c8",x"fd",x"49"),
  3032 => (x"48",x"d0",x"ff",x"87"),
  3033 => (x"f0",x"c3",x"78",x"c4"),
  3034 => (x"66",x"d4",x"1e",x"d2"),
  3035 => (x"de",x"eb",x"fd",x"49"),
  3036 => (x"d8",x"1e",x"c1",x"87"),
  3037 => (x"e8",x"fd",x"49",x"66"),
  3038 => (x"86",x"cc",x"87",x"f1"),
  3039 => (x"c1",x"48",x"66",x"dc"),
  3040 => (x"a6",x"e0",x"c0",x"80"),
  3041 => (x"02",x"ab",x"c1",x"58"),
  3042 => (x"cc",x"87",x"f3",x"c0"),
  3043 => (x"e0",x"c2",x"49",x"66"),
  3044 => (x"48",x"66",x"d0",x"81"),
  3045 => (x"dd",x"05",x"a8",x"69"),
  3046 => (x"48",x"a6",x"d0",x"87"),
  3047 => (x"cc",x"85",x"78",x"c1"),
  3048 => (x"dc",x"c2",x"49",x"66"),
  3049 => (x"05",x"ad",x"69",x"81"),
  3050 => (x"4d",x"c0",x"87",x"d4"),
  3051 => (x"c1",x"48",x"66",x"d4"),
  3052 => (x"58",x"a6",x"d8",x"80"),
  3053 => (x"66",x"d0",x"87",x"c8"),
  3054 => (x"d4",x"80",x"c1",x"48"),
  3055 => (x"8b",x"c1",x"58",x"a6"),
  3056 => (x"eb",x"fd",x"05",x"8c"),
  3057 => (x"02",x"66",x"d8",x"87"),
  3058 => (x"66",x"dc",x"87",x"da"),
  3059 => (x"99",x"ff",x"c3",x"49"),
  3060 => (x"dc",x"59",x"a6",x"d4"),
  3061 => (x"b7",x"c8",x"49",x"66"),
  3062 => (x"59",x"a6",x"d8",x"29"),
  3063 => (x"d8",x"49",x"66",x"dc"),
  3064 => (x"4d",x"71",x"29",x"b7"),
  3065 => (x"49",x"bf",x"97",x"6e"),
  3066 => (x"75",x"99",x"f0",x"c3"),
  3067 => (x"d8",x"1e",x"71",x"b1"),
  3068 => (x"b7",x"c8",x"49",x"66"),
  3069 => (x"dc",x"1e",x"71",x"29"),
  3070 => (x"66",x"dc",x"1e",x"66"),
  3071 => (x"97",x"66",x"d4",x"1e"),
  3072 => (x"c0",x"1e",x"49",x"bf"),
  3073 => (x"87",x"fe",x"e9",x"49"),
  3074 => (x"9b",x"73",x"86",x"d4"),
  3075 => (x"d0",x"87",x"c7",x"02"),
  3076 => (x"87",x"fc",x"e1",x"49"),
  3077 => (x"d0",x"c2",x"87",x"c6"),
  3078 => (x"87",x"f4",x"e1",x"49"),
  3079 => (x"fb",x"05",x"9b",x"73"),
  3080 => (x"8e",x"e0",x"87",x"e1"),
  3081 => (x"0e",x"87",x"cc",x"e7"),
  3082 => (x"5d",x"5c",x"5b",x"5e"),
  3083 => (x"71",x"86",x"f8",x"0e"),
  3084 => (x"49",x"a4",x"c8",x"4c"),
  3085 => (x"2a",x"c9",x"4a",x"69"),
  3086 => (x"c3",x"02",x"9a",x"72"),
  3087 => (x"1e",x"72",x"87",x"ca"),
  3088 => (x"4a",x"d1",x"49",x"72"),
  3089 => (x"87",x"c8",x"c3",x"fd"),
  3090 => (x"99",x"71",x"4a",x"26"),
  3091 => (x"87",x"c4",x"c2",x"05"),
  3092 => (x"c0",x"c0",x"c4",x"c1"),
  3093 => (x"fb",x"c1",x"01",x"aa"),
  3094 => (x"cc",x"7e",x"d1",x"87"),
  3095 => (x"01",x"aa",x"c0",x"f0"),
  3096 => (x"4d",x"c4",x"87",x"c5"),
  3097 => (x"72",x"87",x"cc",x"c1"),
  3098 => (x"c6",x"49",x"72",x"1e"),
  3099 => (x"df",x"c2",x"fd",x"4a"),
  3100 => (x"71",x"4a",x"26",x"87"),
  3101 => (x"87",x"cc",x"05",x"99"),
  3102 => (x"aa",x"c0",x"e0",x"d9"),
  3103 => (x"c6",x"87",x"c5",x"01"),
  3104 => (x"87",x"ef",x"c0",x"4d"),
  3105 => (x"1e",x"72",x"4b",x"c5"),
  3106 => (x"4a",x"73",x"49",x"72"),
  3107 => (x"87",x"c0",x"c2",x"fd"),
  3108 => (x"99",x"71",x"4a",x"26"),
  3109 => (x"73",x"87",x"cb",x"05"),
  3110 => (x"c0",x"d0",x"c4",x"49"),
  3111 => (x"06",x"aa",x"71",x"91"),
  3112 => (x"ab",x"c5",x"87",x"cf"),
  3113 => (x"c1",x"87",x"c2",x"05"),
  3114 => (x"d0",x"83",x"c1",x"83"),
  3115 => (x"d5",x"ff",x"04",x"ab"),
  3116 => (x"72",x"4d",x"73",x"87"),
  3117 => (x"75",x"49",x"72",x"1e"),
  3118 => (x"d3",x"c1",x"fd",x"4a"),
  3119 => (x"26",x"49",x"70",x"87"),
  3120 => (x"72",x"1e",x"71",x"4a"),
  3121 => (x"fd",x"4a",x"d1",x"1e"),
  3122 => (x"26",x"87",x"c5",x"c1"),
  3123 => (x"c8",x"49",x"26",x"4a"),
  3124 => (x"87",x"db",x"58",x"a6"),
  3125 => (x"d0",x"7e",x"ff",x"c0"),
  3126 => (x"c4",x"49",x"72",x"4d"),
  3127 => (x"72",x"1e",x"71",x"29"),
  3128 => (x"4a",x"ff",x"c0",x"1e"),
  3129 => (x"87",x"e8",x"c0",x"fd"),
  3130 => (x"49",x"26",x"4a",x"26"),
  3131 => (x"c2",x"58",x"a6",x"c8"),
  3132 => (x"c4",x"49",x"a4",x"d8"),
  3133 => (x"dc",x"c2",x"79",x"66"),
  3134 => (x"79",x"75",x"49",x"a4"),
  3135 => (x"49",x"a4",x"e0",x"c2"),
  3136 => (x"e4",x"c2",x"79",x"6e"),
  3137 => (x"79",x"c1",x"49",x"a4"),
  3138 => (x"e6",x"e3",x"8e",x"f8"),
  3139 => (x"49",x"c0",x"1e",x"87"),
  3140 => (x"bf",x"da",x"c6",x"c4"),
  3141 => (x"c1",x"87",x"c2",x"02"),
  3142 => (x"c2",x"c9",x"c4",x"49"),
  3143 => (x"87",x"c2",x"02",x"bf"),
  3144 => (x"d0",x"ff",x"b1",x"c2"),
  3145 => (x"78",x"c5",x"c8",x"48"),
  3146 => (x"c3",x"48",x"d4",x"ff"),
  3147 => (x"78",x"71",x"78",x"fa"),
  3148 => (x"c4",x"48",x"d0",x"ff"),
  3149 => (x"1e",x"4f",x"26",x"78"),
  3150 => (x"4a",x"71",x"1e",x"73"),
  3151 => (x"49",x"66",x"cc",x"1e"),
  3152 => (x"c4",x"91",x"e8",x"c2"),
  3153 => (x"71",x"4b",x"d2",x"c6"),
  3154 => (x"fd",x"49",x"73",x"83"),
  3155 => (x"c4",x"87",x"f0",x"de"),
  3156 => (x"02",x"98",x"70",x"86"),
  3157 => (x"49",x"73",x"87",x"cb"),
  3158 => (x"87",x"f5",x"e7",x"fd"),
  3159 => (x"c6",x"fb",x"49",x"73"),
  3160 => (x"87",x"e9",x"fe",x"87"),
  3161 => (x"0e",x"87",x"d0",x"e2"),
  3162 => (x"5d",x"5c",x"5b",x"5e"),
  3163 => (x"ff",x"86",x"f4",x"0e"),
  3164 => (x"70",x"87",x"f5",x"dc"),
  3165 => (x"02",x"99",x"c4",x"49"),
  3166 => (x"ff",x"87",x"ec",x"c5"),
  3167 => (x"c5",x"c8",x"48",x"d0"),
  3168 => (x"48",x"d4",x"ff",x"78"),
  3169 => (x"c0",x"78",x"c0",x"c2"),
  3170 => (x"78",x"78",x"78",x"78"),
  3171 => (x"d4",x"ff",x"4d",x"78"),
  3172 => (x"76",x"78",x"c0",x"48"),
  3173 => (x"ff",x"49",x"a5",x"4a"),
  3174 => (x"79",x"97",x"bf",x"d4"),
  3175 => (x"c0",x"48",x"d4",x"ff"),
  3176 => (x"c1",x"51",x"68",x"78"),
  3177 => (x"ad",x"b7",x"c8",x"85"),
  3178 => (x"ff",x"87",x"e3",x"04"),
  3179 => (x"78",x"c4",x"48",x"d0"),
  3180 => (x"48",x"66",x"97",x"c6"),
  3181 => (x"70",x"58",x"a6",x"cc"),
  3182 => (x"c4",x"9b",x"d0",x"4b"),
  3183 => (x"49",x"73",x"2b",x"b7"),
  3184 => (x"c4",x"91",x"e8",x"c2"),
  3185 => (x"c8",x"81",x"d2",x"c6"),
  3186 => (x"ca",x"05",x"69",x"81"),
  3187 => (x"49",x"d1",x"c2",x"87"),
  3188 => (x"87",x"fc",x"da",x"ff"),
  3189 => (x"c7",x"87",x"d0",x"c4"),
  3190 => (x"49",x"4c",x"66",x"97"),
  3191 => (x"d0",x"99",x"f0",x"c3"),
  3192 => (x"87",x"cc",x"05",x"a9"),
  3193 => (x"49",x"72",x"1e",x"73"),
  3194 => (x"c4",x"87",x"d2",x"e3"),
  3195 => (x"87",x"f7",x"c3",x"86"),
  3196 => (x"05",x"ac",x"d0",x"c2"),
  3197 => (x"49",x"72",x"87",x"c8"),
  3198 => (x"c3",x"87",x"e5",x"e3"),
  3199 => (x"ec",x"c3",x"87",x"e9"),
  3200 => (x"87",x"ce",x"05",x"ac"),
  3201 => (x"1e",x"73",x"1e",x"c0"),
  3202 => (x"cf",x"e4",x"49",x"72"),
  3203 => (x"c3",x"86",x"c8",x"87"),
  3204 => (x"d1",x"c2",x"87",x"d5"),
  3205 => (x"87",x"cc",x"05",x"ac"),
  3206 => (x"49",x"72",x"1e",x"73"),
  3207 => (x"c4",x"87",x"e9",x"e5"),
  3208 => (x"87",x"c3",x"c3",x"86"),
  3209 => (x"05",x"ac",x"c6",x"c3"),
  3210 => (x"1e",x"73",x"87",x"cc"),
  3211 => (x"cc",x"e6",x"49",x"72"),
  3212 => (x"c2",x"86",x"c4",x"87"),
  3213 => (x"e0",x"c0",x"87",x"f1"),
  3214 => (x"87",x"cf",x"05",x"ac"),
  3215 => (x"73",x"1e",x"1e",x"c0"),
  3216 => (x"e8",x"49",x"72",x"1e"),
  3217 => (x"86",x"cc",x"87",x"f3"),
  3218 => (x"c3",x"87",x"dc",x"c2"),
  3219 => (x"d0",x"05",x"ac",x"c4"),
  3220 => (x"c1",x"1e",x"c0",x"87"),
  3221 => (x"72",x"1e",x"73",x"1e"),
  3222 => (x"87",x"dd",x"e8",x"49"),
  3223 => (x"c6",x"c2",x"86",x"cc"),
  3224 => (x"ac",x"f0",x"c0",x"87"),
  3225 => (x"c0",x"87",x"ce",x"05"),
  3226 => (x"72",x"1e",x"73",x"1e"),
  3227 => (x"87",x"c2",x"f0",x"49"),
  3228 => (x"f2",x"c1",x"86",x"c8"),
  3229 => (x"ac",x"c5",x"c3",x"87"),
  3230 => (x"c1",x"87",x"ce",x"05"),
  3231 => (x"72",x"1e",x"73",x"1e"),
  3232 => (x"87",x"ee",x"ef",x"49"),
  3233 => (x"de",x"c1",x"86",x"c8"),
  3234 => (x"05",x"ac",x"c8",x"87"),
  3235 => (x"1e",x"73",x"87",x"cc"),
  3236 => (x"d3",x"e6",x"49",x"72"),
  3237 => (x"c1",x"86",x"c4",x"87"),
  3238 => (x"c0",x"c1",x"87",x"cd"),
  3239 => (x"87",x"d0",x"05",x"ac"),
  3240 => (x"1e",x"c0",x"1e",x"c1"),
  3241 => (x"49",x"72",x"1e",x"73"),
  3242 => (x"cc",x"87",x"ce",x"e7"),
  3243 => (x"87",x"f7",x"c0",x"86"),
  3244 => (x"cc",x"05",x"9c",x"74"),
  3245 => (x"72",x"1e",x"73",x"87"),
  3246 => (x"87",x"f1",x"e4",x"49"),
  3247 => (x"e6",x"c0",x"86",x"c4"),
  3248 => (x"1e",x"66",x"c8",x"87"),
  3249 => (x"49",x"66",x"97",x"c9"),
  3250 => (x"66",x"97",x"cc",x"1e"),
  3251 => (x"97",x"cf",x"1e",x"49"),
  3252 => (x"d2",x"1e",x"49",x"66"),
  3253 => (x"1e",x"49",x"66",x"97"),
  3254 => (x"de",x"ff",x"49",x"c4"),
  3255 => (x"86",x"d4",x"87",x"e8"),
  3256 => (x"ff",x"49",x"d1",x"c2"),
  3257 => (x"f4",x"87",x"e9",x"d6"),
  3258 => (x"c6",x"dc",x"ff",x"8e"),
  3259 => (x"5b",x"5e",x"0e",x"87"),
  3260 => (x"1e",x"0e",x"5d",x"5c"),
  3261 => (x"d4",x"ff",x"7e",x"71"),
  3262 => (x"c4",x"1e",x"6e",x"4b"),
  3263 => (x"fd",x"49",x"e2",x"cb"),
  3264 => (x"c4",x"87",x"fc",x"d7"),
  3265 => (x"9d",x"4d",x"70",x"86"),
  3266 => (x"87",x"c3",x"c3",x"02"),
  3267 => (x"bf",x"ea",x"cb",x"c4"),
  3268 => (x"fd",x"49",x"6e",x"4c"),
  3269 => (x"ff",x"87",x"cf",x"f4"),
  3270 => (x"c5",x"c8",x"48",x"d0"),
  3271 => (x"7b",x"d6",x"c1",x"78"),
  3272 => (x"7b",x"15",x"4a",x"c0"),
  3273 => (x"e0",x"c0",x"82",x"c1"),
  3274 => (x"f5",x"04",x"aa",x"b7"),
  3275 => (x"48",x"d0",x"ff",x"87"),
  3276 => (x"c5",x"c8",x"78",x"c4"),
  3277 => (x"7b",x"d3",x"c1",x"78"),
  3278 => (x"78",x"c4",x"7b",x"c1"),
  3279 => (x"c1",x"02",x"9c",x"74"),
  3280 => (x"f0",x"c3",x"87",x"fc"),
  3281 => (x"c0",x"c8",x"7e",x"d2"),
  3282 => (x"b7",x"c0",x"8c",x"4d"),
  3283 => (x"87",x"c6",x"03",x"ac"),
  3284 => (x"4d",x"a4",x"c0",x"c8"),
  3285 => (x"fd",x"c3",x"4c",x"c0"),
  3286 => (x"49",x"bf",x"97",x"c3"),
  3287 => (x"d2",x"02",x"99",x"d0"),
  3288 => (x"c4",x"1e",x"c0",x"87"),
  3289 => (x"fd",x"49",x"e2",x"cb"),
  3290 => (x"c4",x"87",x"e1",x"da"),
  3291 => (x"4a",x"49",x"70",x"86"),
  3292 => (x"c3",x"87",x"ef",x"c0"),
  3293 => (x"c4",x"1e",x"d2",x"f0"),
  3294 => (x"fd",x"49",x"e2",x"cb"),
  3295 => (x"c4",x"87",x"cd",x"da"),
  3296 => (x"4a",x"49",x"70",x"86"),
  3297 => (x"c8",x"48",x"d0",x"ff"),
  3298 => (x"d4",x"c1",x"78",x"c5"),
  3299 => (x"bf",x"97",x"6e",x"7b"),
  3300 => (x"c1",x"48",x"6e",x"7b"),
  3301 => (x"c1",x"7e",x"70",x"80"),
  3302 => (x"f0",x"ff",x"05",x"8d"),
  3303 => (x"48",x"d0",x"ff",x"87"),
  3304 => (x"9a",x"72",x"78",x"c4"),
  3305 => (x"c0",x"87",x"c5",x"05"),
  3306 => (x"87",x"e5",x"c0",x"48"),
  3307 => (x"cb",x"c4",x"1e",x"c1"),
  3308 => (x"d7",x"fd",x"49",x"e2"),
  3309 => (x"86",x"c4",x"87",x"f5"),
  3310 => (x"fe",x"05",x"9c",x"74"),
  3311 => (x"d0",x"ff",x"87",x"c4"),
  3312 => (x"78",x"c5",x"c8",x"48"),
  3313 => (x"c0",x"7b",x"d3",x"c1"),
  3314 => (x"c1",x"78",x"c4",x"7b"),
  3315 => (x"c0",x"87",x"c2",x"48"),
  3316 => (x"4d",x"26",x"26",x"48"),
  3317 => (x"4b",x"26",x"4c",x"26"),
  3318 => (x"1e",x"00",x"4f",x"26"),
  3319 => (x"bf",x"c4",x"d0",x"c3"),
  3320 => (x"c3",x"b9",x"c1",x"49"),
  3321 => (x"ff",x"59",x"c8",x"d0"),
  3322 => (x"ff",x"c3",x"48",x"d4"),
  3323 => (x"48",x"d0",x"ff",x"78"),
  3324 => (x"ff",x"78",x"e1",x"c8"),
  3325 => (x"78",x"c1",x"48",x"d4"),
  3326 => (x"78",x"71",x"31",x"c4"),
  3327 => (x"c0",x"48",x"d0",x"ff"),
  3328 => (x"4f",x"26",x"78",x"e0"),
  3329 => (x"00",x"00",x"00",x"00"),
  3330 => (x"5c",x"5b",x"5e",x"0e"),
  3331 => (x"4c",x"71",x"1e",x"0e"),
  3332 => (x"87",x"cc",x"fd",x"fe"),
  3333 => (x"66",x"d0",x"4b",x"70"),
  3334 => (x"ef",x"c0",x"c4",x"1e"),
  3335 => (x"e2",x"dc",x"fe",x"49"),
  3336 => (x"73",x"86",x"c4",x"87"),
  3337 => (x"87",x"d9",x"05",x"9b"),
  3338 => (x"4a",x"a4",x"f4",x"c0"),
  3339 => (x"49",x"a4",x"f0",x"c0"),
  3340 => (x"66",x"d0",x"82",x"69"),
  3341 => (x"c1",x"48",x"69",x"52"),
  3342 => (x"6e",x"7e",x"70",x"80"),
  3343 => (x"70",x"98",x"cf",x"48"),
  3344 => (x"87",x"c2",x"26",x"79"),
  3345 => (x"4c",x"26",x"4d",x"26"),
  3346 => (x"4f",x"26",x"4b",x"26"),
  3347 => (x"5c",x"5b",x"5e",x"0e"),
  3348 => (x"cc",x"4b",x"71",x"0e"),
  3349 => (x"c2",x"49",x"4c",x"66"),
  3350 => (x"ca",x"02",x"99",x"c0"),
  3351 => (x"1e",x"e0",x"c3",x"87"),
  3352 => (x"e3",x"fe",x"49",x"73"),
  3353 => (x"74",x"86",x"c4",x"87"),
  3354 => (x"99",x"c0",x"c4",x"49"),
  3355 => (x"c2",x"87",x"c5",x"02"),
  3356 => (x"87",x"c3",x"b4",x"c0"),
  3357 => (x"74",x"9c",x"ff",x"c1"),
  3358 => (x"fe",x"49",x"73",x"1e"),
  3359 => (x"ff",x"26",x"87",x"ca"),
  3360 => (x"73",x"1e",x"87",x"c4"),
  3361 => (x"d3",x"c3",x"1e",x"1e"),
  3362 => (x"ff",x"49",x"bf",x"e8"),
  3363 => (x"70",x"87",x"c8",x"c8"),
  3364 => (x"cf",x"c1",x"02",x"98"),
  3365 => (x"e6",x"ce",x"c4",x"87"),
  3366 => (x"ce",x"c4",x"48",x"bf"),
  3367 => (x"02",x"a8",x"bf",x"ea"),
  3368 => (x"c4",x"87",x"c1",x"c1"),
  3369 => (x"c4",x"4b",x"ee",x"ce"),
  3370 => (x"83",x"bf",x"e6",x"ce"),
  3371 => (x"c0",x"4b",x"6b",x"97"),
  3372 => (x"c7",x"ff",x"49",x"e8"),
  3373 => (x"49",x"70",x"87",x"d5"),
  3374 => (x"59",x"ec",x"d3",x"c3"),
  3375 => (x"c8",x"48",x"d0",x"ff"),
  3376 => (x"d4",x"ff",x"78",x"e1"),
  3377 => (x"73",x"78",x"c5",x"48"),
  3378 => (x"08",x"d4",x"ff",x"48"),
  3379 => (x"48",x"d0",x"ff",x"78"),
  3380 => (x"c4",x"78",x"e0",x"c0"),
  3381 => (x"48",x"bf",x"e6",x"ce"),
  3382 => (x"7e",x"70",x"80",x"c1"),
  3383 => (x"98",x"cf",x"48",x"6e"),
  3384 => (x"58",x"ea",x"ce",x"c4"),
  3385 => (x"87",x"e0",x"fd",x"26"),
  3386 => (x"00",x"00",x"00",x"00"),
  3387 => (x"5c",x"5b",x"5e",x"0e"),
  3388 => (x"d8",x"ff",x"0e",x"5d"),
  3389 => (x"c4",x"7e",x"c0",x"86"),
  3390 => (x"49",x"bf",x"fe",x"cd"),
  3391 => (x"1e",x"71",x"81",x"c2"),
  3392 => (x"4a",x"c6",x"1e",x"72"),
  3393 => (x"87",x"fc",x"f0",x"fc"),
  3394 => (x"4a",x"26",x"48",x"71"),
  3395 => (x"a6",x"c8",x"49",x"26"),
  3396 => (x"fe",x"cd",x"c4",x"58"),
  3397 => (x"81",x"c4",x"49",x"bf"),
  3398 => (x"1e",x"72",x"1e",x"71"),
  3399 => (x"f0",x"fc",x"4a",x"c6"),
  3400 => (x"48",x"71",x"87",x"e2"),
  3401 => (x"49",x"26",x"4a",x"26"),
  3402 => (x"fd",x"58",x"a6",x"cc"),
  3403 => (x"df",x"c3",x"87",x"d4"),
  3404 => (x"ff",x"49",x"bf",x"f6"),
  3405 => (x"70",x"87",x"e0",x"c5"),
  3406 => (x"f3",x"ca",x"02",x"98"),
  3407 => (x"ff",x"49",x"d0",x"87"),
  3408 => (x"70",x"87",x"c8",x"c5"),
  3409 => (x"fa",x"df",x"c3",x"49"),
  3410 => (x"74",x"4c",x"c0",x"59"),
  3411 => (x"fe",x"91",x"c4",x"49"),
  3412 => (x"4a",x"69",x"81",x"d0"),
  3413 => (x"cd",x"c4",x"49",x"74"),
  3414 => (x"c4",x"81",x"bf",x"fe"),
  3415 => (x"ce",x"ce",x"c4",x"91"),
  3416 => (x"9a",x"79",x"72",x"81"),
  3417 => (x"72",x"87",x"d2",x"02"),
  3418 => (x"71",x"89",x"c1",x"49"),
  3419 => (x"c1",x"48",x"6e",x"9a"),
  3420 => (x"72",x"7e",x"70",x"80"),
  3421 => (x"ee",x"ff",x"05",x"9a"),
  3422 => (x"c2",x"84",x"c1",x"87"),
  3423 => (x"ff",x"04",x"ac",x"b7"),
  3424 => (x"48",x"6e",x"87",x"c9"),
  3425 => (x"a8",x"b7",x"fc",x"c0"),
  3426 => (x"87",x"e4",x"c9",x"04"),
  3427 => (x"4a",x"74",x"4c",x"c0"),
  3428 => (x"c4",x"82",x"66",x"c4"),
  3429 => (x"ce",x"ce",x"c4",x"92"),
  3430 => (x"c8",x"49",x"74",x"82"),
  3431 => (x"91",x"c4",x"81",x"66"),
  3432 => (x"81",x"ce",x"ce",x"c4"),
  3433 => (x"49",x"69",x"4a",x"6a"),
  3434 => (x"4b",x"74",x"b9",x"72"),
  3435 => (x"bf",x"fe",x"cd",x"c4"),
  3436 => (x"c4",x"93",x"c4",x"83"),
  3437 => (x"6b",x"83",x"ce",x"ce"),
  3438 => (x"71",x"48",x"72",x"ba"),
  3439 => (x"58",x"a6",x"d4",x"98"),
  3440 => (x"cd",x"c4",x"49",x"74"),
  3441 => (x"c4",x"81",x"bf",x"fe"),
  3442 => (x"ce",x"ce",x"c4",x"91"),
  3443 => (x"d4",x"7e",x"69",x"81"),
  3444 => (x"78",x"c0",x"48",x"a6"),
  3445 => (x"c3",x"5c",x"a6",x"d0"),
  3446 => (x"66",x"d0",x"4c",x"ff"),
  3447 => (x"02",x"29",x"df",x"49"),
  3448 => (x"cc",x"87",x"dc",x"c7"),
  3449 => (x"e0",x"c0",x"4a",x"66"),
  3450 => (x"82",x"66",x"d4",x"92"),
  3451 => (x"72",x"48",x"ff",x"c0"),
  3452 => (x"d8",x"4a",x"70",x"88"),
  3453 => (x"78",x"c0",x"48",x"a6"),
  3454 => (x"78",x"c0",x"80",x"c4"),
  3455 => (x"29",x"df",x"49",x"6e"),
  3456 => (x"59",x"a6",x"e4",x"c0"),
  3457 => (x"48",x"fa",x"cd",x"c4"),
  3458 => (x"49",x"72",x"78",x"c1"),
  3459 => (x"2a",x"b7",x"31",x"c3"),
  3460 => (x"ff",x"c0",x"b1",x"72"),
  3461 => (x"c3",x"91",x"c4",x"99"),
  3462 => (x"71",x"4d",x"ec",x"eb"),
  3463 => (x"49",x"4b",x"6d",x"85"),
  3464 => (x"99",x"c0",x"c0",x"c4"),
  3465 => (x"c0",x"87",x"d7",x"02"),
  3466 => (x"c0",x"02",x"66",x"e0"),
  3467 => (x"80",x"c8",x"87",x"c7"),
  3468 => (x"ca",x"c6",x"78",x"c0"),
  3469 => (x"c2",x"ce",x"c4",x"87"),
  3470 => (x"c6",x"78",x"c1",x"48"),
  3471 => (x"e0",x"c0",x"87",x"c1"),
  3472 => (x"87",x"d8",x"02",x"66"),
  3473 => (x"c0",x"c2",x"49",x"73"),
  3474 => (x"c0",x"02",x"99",x"c0"),
  3475 => (x"b7",x"d0",x"87",x"c3"),
  3476 => (x"fd",x"48",x"6d",x"2b"),
  3477 => (x"70",x"98",x"ff",x"ff"),
  3478 => (x"87",x"fa",x"c0",x"7d"),
  3479 => (x"bf",x"c2",x"ce",x"c4"),
  3480 => (x"87",x"f2",x"c0",x"02"),
  3481 => (x"b7",x"d0",x"48",x"73"),
  3482 => (x"a6",x"e8",x"c0",x"28"),
  3483 => (x"02",x"98",x"70",x"58"),
  3484 => (x"c4",x"87",x"e3",x"c0"),
  3485 => (x"49",x"bf",x"ca",x"ce"),
  3486 => (x"99",x"c0",x"e0",x"c0"),
  3487 => (x"87",x"ca",x"c0",x"02"),
  3488 => (x"e0",x"c0",x"49",x"70"),
  3489 => (x"c0",x"02",x"99",x"c0"),
  3490 => (x"48",x"6d",x"87",x"cc"),
  3491 => (x"b0",x"c0",x"c0",x"c2"),
  3492 => (x"e4",x"c0",x"7d",x"70"),
  3493 => (x"49",x"73",x"4b",x"66"),
  3494 => (x"99",x"c0",x"c0",x"c8"),
  3495 => (x"87",x"ff",x"c2",x"02"),
  3496 => (x"02",x"66",x"e0",x"c0"),
  3497 => (x"73",x"87",x"c8",x"c0"),
  3498 => (x"9a",x"c0",x"cc",x"4a"),
  3499 => (x"f3",x"87",x"cf",x"c0"),
  3500 => (x"ce",x"c4",x"9b",x"ff"),
  3501 => (x"cc",x"4a",x"bf",x"ca"),
  3502 => (x"b3",x"72",x"9a",x"c0"),
  3503 => (x"9a",x"72",x"7d",x"73"),
  3504 => (x"48",x"87",x"df",x"02"),
  3505 => (x"c0",x"88",x"c0",x"c4"),
  3506 => (x"70",x"58",x"a6",x"e8"),
  3507 => (x"e0",x"c0",x"02",x"98"),
  3508 => (x"c0",x"c4",x"48",x"87"),
  3509 => (x"a6",x"e8",x"c0",x"88"),
  3510 => (x"02",x"98",x"70",x"58"),
  3511 => (x"c1",x"87",x"c2",x"c1"),
  3512 => (x"49",x"73",x"87",x"ef"),
  3513 => (x"91",x"c2",x"99",x"74"),
  3514 => (x"81",x"e0",x"eb",x"c3"),
  3515 => (x"ee",x"c1",x"4b",x"11"),
  3516 => (x"74",x"49",x"73",x"87"),
  3517 => (x"c3",x"91",x"c2",x"99"),
  3518 => (x"c1",x"81",x"e0",x"eb"),
  3519 => (x"c4",x"4b",x"11",x"81"),
  3520 => (x"49",x"bf",x"ca",x"ce"),
  3521 => (x"c0",x"99",x"c0",x"c4"),
  3522 => (x"02",x"99",x"66",x"e0"),
  3523 => (x"dc",x"87",x"c9",x"c0"),
  3524 => (x"ea",x"c0",x"48",x"a6"),
  3525 => (x"87",x"c7",x"c1",x"78"),
  3526 => (x"c4",x"48",x"a6",x"d8"),
  3527 => (x"fe",x"c0",x"78",x"ea"),
  3528 => (x"74",x"49",x"73",x"87"),
  3529 => (x"c3",x"91",x"c2",x"99"),
  3530 => (x"c1",x"81",x"e0",x"eb"),
  3531 => (x"c4",x"4b",x"11",x"81"),
  3532 => (x"49",x"bf",x"ca",x"ce"),
  3533 => (x"c0",x"99",x"c0",x"c8"),
  3534 => (x"02",x"99",x"66",x"e0"),
  3535 => (x"dc",x"87",x"c9",x"c0"),
  3536 => (x"f6",x"c0",x"48",x"a6"),
  3537 => (x"87",x"d7",x"c0",x"78"),
  3538 => (x"c4",x"48",x"a6",x"d8"),
  3539 => (x"ce",x"c0",x"78",x"f6"),
  3540 => (x"74",x"49",x"73",x"87"),
  3541 => (x"c3",x"91",x"c2",x"99"),
  3542 => (x"c1",x"81",x"e0",x"eb"),
  3543 => (x"c0",x"4b",x"11",x"81"),
  3544 => (x"c0",x"02",x"66",x"e0"),
  3545 => (x"49",x"73",x"87",x"db"),
  3546 => (x"fc",x"c7",x"b9",x"ff"),
  3547 => (x"48",x"71",x"99",x"c0"),
  3548 => (x"bf",x"ca",x"ce",x"c4"),
  3549 => (x"ce",x"ce",x"c4",x"98"),
  3550 => (x"c4",x"9b",x"74",x"58"),
  3551 => (x"d3",x"c0",x"b3",x"c0"),
  3552 => (x"c7",x"49",x"73",x"87"),
  3553 => (x"71",x"99",x"c0",x"fc"),
  3554 => (x"ca",x"ce",x"c4",x"48"),
  3555 => (x"ce",x"c4",x"b0",x"bf"),
  3556 => (x"9b",x"74",x"58",x"ce"),
  3557 => (x"c0",x"02",x"66",x"d8"),
  3558 => (x"c4",x"1e",x"87",x"ca"),
  3559 => (x"f2",x"49",x"fa",x"cd"),
  3560 => (x"86",x"c4",x"87",x"ea"),
  3561 => (x"cd",x"c4",x"1e",x"73"),
  3562 => (x"df",x"f2",x"49",x"fa"),
  3563 => (x"dc",x"86",x"c4",x"87"),
  3564 => (x"ca",x"c0",x"02",x"66"),
  3565 => (x"cd",x"c4",x"1e",x"87"),
  3566 => (x"cf",x"f2",x"49",x"fa"),
  3567 => (x"d0",x"86",x"c4",x"87"),
  3568 => (x"30",x"c1",x"48",x"66"),
  3569 => (x"6e",x"58",x"a6",x"d4"),
  3570 => (x"70",x"30",x"c1",x"48"),
  3571 => (x"48",x"66",x"d4",x"7e"),
  3572 => (x"a6",x"d8",x"80",x"c1"),
  3573 => (x"b7",x"e0",x"c0",x"58"),
  3574 => (x"fd",x"f7",x"04",x"a8"),
  3575 => (x"4c",x"66",x"cc",x"87"),
  3576 => (x"b7",x"c2",x"84",x"c1"),
  3577 => (x"e5",x"f6",x"04",x"ac"),
  3578 => (x"fe",x"cd",x"c4",x"87"),
  3579 => (x"78",x"66",x"c4",x"48"),
  3580 => (x"f1",x"8e",x"d8",x"ff"),
  3581 => (x"00",x"00",x"87",x"ce"),
  3582 => (x"c0",x"1e",x"00",x"00"),
  3583 => (x"c4",x"49",x"72",x"4a"),
  3584 => (x"ce",x"ce",x"c4",x"91"),
  3585 => (x"c1",x"79",x"ff",x"81"),
  3586 => (x"aa",x"b7",x"c6",x"82"),
  3587 => (x"c4",x"87",x"ee",x"04"),
  3588 => (x"c0",x"48",x"fe",x"cd"),
  3589 => (x"80",x"c8",x"78",x"40"),
  3590 => (x"4f",x"26",x"78",x"c0"),
  3591 => (x"71",x"1e",x"73",x"1e"),
  3592 => (x"87",x"c8",x"f3",x"4b"),
  3593 => (x"d0",x"fe",x"49",x"73"),
  3594 => (x"db",x"f0",x"87",x"ca"),
  3595 => (x"5b",x"5e",x"0e",x"87"),
  3596 => (x"71",x"1e",x"0e",x"5c"),
  3597 => (x"d0",x"4b",x"c0",x"4c"),
  3598 => (x"e9",x"c0",x"02",x"66"),
  3599 => (x"8a",x"c1",x"4a",x"87"),
  3600 => (x"87",x"e2",x"c0",x"02"),
  3601 => (x"87",x"de",x"02",x"8a"),
  3602 => (x"02",x"8a",x"ee",x"c0"),
  3603 => (x"c1",x"87",x"c6",x"c1"),
  3604 => (x"72",x"7e",x"73",x"8a"),
  3605 => (x"d7",x"c1",x"02",x"9a"),
  3606 => (x"73",x"8a",x"c1",x"87"),
  3607 => (x"02",x"9a",x"72",x"7e"),
  3608 => (x"c1",x"87",x"cd",x"c1"),
  3609 => (x"9c",x"74",x"87",x"d9"),
  3610 => (x"87",x"d3",x"c1",x"02"),
  3611 => (x"c1",x"02",x"6c",x"97"),
  3612 => (x"c0",x"c4",x"87",x"cd"),
  3613 => (x"c1",x"48",x"bf",x"f9"),
  3614 => (x"fd",x"c0",x"c4",x"b0"),
  3615 => (x"c0",x"d6",x"fe",x"58"),
  3616 => (x"49",x"66",x"d0",x"87"),
  3617 => (x"cf",x"c3",x"81",x"c1"),
  3618 => (x"74",x"59",x"97",x"de"),
  3619 => (x"87",x"dd",x"e9",x"49"),
  3620 => (x"ea",x"c0",x"4b",x"70"),
  3621 => (x"4b",x"66",x"d0",x"87"),
  3622 => (x"73",x"8b",x"f0",x"c0"),
  3623 => (x"fe",x"49",x"c0",x"1e"),
  3624 => (x"73",x"87",x"eb",x"fd"),
  3625 => (x"fe",x"49",x"74",x"1e"),
  3626 => (x"c8",x"87",x"e3",x"fd"),
  3627 => (x"87",x"e0",x"c0",x"86"),
  3628 => (x"c0",x"49",x"66",x"d0"),
  3629 => (x"1e",x"71",x"89",x"f1"),
  3630 => (x"fa",x"e1",x"49",x"74"),
  3631 => (x"c4",x"86",x"c4",x"87"),
  3632 => (x"48",x"bf",x"f9",x"c0"),
  3633 => (x"c0",x"c4",x"98",x"fe"),
  3634 => (x"d4",x"fe",x"58",x"fd"),
  3635 => (x"48",x"73",x"87",x"f3"),
  3636 => (x"87",x"f2",x"ed",x"26"),
  3637 => (x"c0",x"1e",x"73",x"1e"),
  3638 => (x"f9",x"c0",x"c4",x"4b"),
  3639 => (x"b0",x"c1",x"48",x"bf"),
  3640 => (x"58",x"fd",x"c0",x"c4"),
  3641 => (x"87",x"d9",x"d4",x"fe"),
  3642 => (x"48",x"cc",x"c4",x"c1"),
  3643 => (x"1e",x"c8",x"50",x"c0"),
  3644 => (x"49",x"fe",x"ce",x"c4"),
  3645 => (x"87",x"ed",x"db",x"fd"),
  3646 => (x"1e",x"72",x"86",x"c4"),
  3647 => (x"48",x"dc",x"e6",x"c3"),
  3648 => (x"49",x"c6",x"cf",x"c4"),
  3649 => (x"20",x"4a",x"a1",x"c4"),
  3650 => (x"05",x"aa",x"71",x"41"),
  3651 => (x"4a",x"26",x"87",x"f9"),
  3652 => (x"49",x"fe",x"ce",x"c4"),
  3653 => (x"87",x"c6",x"fe",x"fc"),
  3654 => (x"02",x"9a",x"4a",x"70"),
  3655 => (x"fd",x"49",x"87",x"c5"),
  3656 => (x"72",x"87",x"f5",x"ce"),
  3657 => (x"e0",x"e6",x"c3",x"1e"),
  3658 => (x"c6",x"cf",x"c4",x"48"),
  3659 => (x"4a",x"a1",x"c4",x"49"),
  3660 => (x"aa",x"71",x"41",x"20"),
  3661 => (x"87",x"f8",x"ff",x"05"),
  3662 => (x"1e",x"c0",x"4a",x"26"),
  3663 => (x"49",x"fe",x"ce",x"c4"),
  3664 => (x"87",x"ca",x"fb",x"fe"),
  3665 => (x"1e",x"72",x"86",x"c4"),
  3666 => (x"48",x"e4",x"e6",x"c3"),
  3667 => (x"49",x"c6",x"cf",x"c4"),
  3668 => (x"20",x"4a",x"a1",x"c4"),
  3669 => (x"05",x"aa",x"71",x"41"),
  3670 => (x"26",x"87",x"f8",x"ff"),
  3671 => (x"fe",x"ce",x"c4",x"4a"),
  3672 => (x"87",x"c9",x"e6",x"49"),
  3673 => (x"c0",x"05",x"98",x"70"),
  3674 => (x"e6",x"c3",x"87",x"c4"),
  3675 => (x"49",x"c0",x"4b",x"e8"),
  3676 => (x"87",x"c6",x"cc",x"fd"),
  3677 => (x"73",x"87",x"c3",x"fa"),
  3678 => (x"c5",x"c0",x"02",x"9b"),
  3679 => (x"db",x"fc",x"49",x"87"),
  3680 => (x"49",x"ca",x"87",x"e7"),
  3681 => (x"87",x"c7",x"db",x"fc"),
  3682 => (x"bf",x"f9",x"c0",x"c4"),
  3683 => (x"c4",x"98",x"fe",x"48"),
  3684 => (x"fe",x"58",x"fd",x"c0"),
  3685 => (x"73",x"87",x"ea",x"d1"),
  3686 => (x"87",x"ec",x"ea",x"48"),
  3687 => (x"00",x"20",x"20",x"20"),
  3688 => (x"00",x"44",x"48",x"56"),
  3689 => (x"00",x"4d",x"4f",x"52"),
  3690 => (x"20",x"4d",x"4f",x"52"),
  3691 => (x"64",x"61",x"6f",x"6c"),
  3692 => (x"20",x"67",x"6e",x"69"),
  3693 => (x"6c",x"69",x"61",x"66"),
  3694 => (x"0e",x"00",x"64",x"65"),
  3695 => (x"5d",x"5c",x"5b",x"5e"),
  3696 => (x"d7",x"c1",x"1e",x"0e"),
  3697 => (x"87",x"f2",x"f8",x"4d"),
  3698 => (x"fe",x"87",x"e1",x"ec"),
  3699 => (x"fe",x"87",x"e9",x"e9"),
  3700 => (x"ff",x"87",x"d1",x"f5"),
  3701 => (x"6e",x"87",x"d0",x"de"),
  3702 => (x"ff",x"ff",x"c1",x"49"),
  3703 => (x"c1",x"48",x"6e",x"99"),
  3704 => (x"71",x"7e",x"70",x"80"),
  3705 => (x"87",x"ca",x"05",x"99"),
  3706 => (x"87",x"e9",x"fd",x"fd"),
  3707 => (x"cf",x"fe",x"49",x"70"),
  3708 => (x"49",x"75",x"87",x"e3"),
  3709 => (x"87",x"c2",x"cc",x"fe"),
  3710 => (x"c2",x"4b",x"49",x"70"),
  3711 => (x"fe",x"49",x"dd",x"9b"),
  3712 => (x"70",x"87",x"f7",x"cb"),
  3713 => (x"ff",x"fe",x"02",x"98"),
  3714 => (x"02",x"9b",x"73",x"87"),
  3715 => (x"75",x"87",x"f9",x"fe"),
  3716 => (x"e5",x"cb",x"fe",x"49"),
  3717 => (x"05",x"98",x"70",x"87"),
  3718 => (x"49",x"dd",x"87",x"cb"),
  3719 => (x"87",x"da",x"cb",x"fe"),
  3720 => (x"de",x"02",x"98",x"70"),
  3721 => (x"fe",x"49",x"c1",x"87"),
  3722 => (x"75",x"87",x"c9",x"c8"),
  3723 => (x"c9",x"cb",x"fe",x"49"),
  3724 => (x"05",x"98",x"70",x"87"),
  3725 => (x"dd",x"87",x"ee",x"ff"),
  3726 => (x"fd",x"ca",x"fe",x"49"),
  3727 => (x"05",x"98",x"70",x"87"),
  3728 => (x"cf",x"87",x"e2",x"ff"),
  3729 => (x"f1",x"fe",x"49",x"e8"),
  3730 => (x"4b",x"70",x"87",x"c1"),
  3731 => (x"eb",x"c3",x"1e",x"c0"),
  3732 => (x"ef",x"fe",x"49",x"c9"),
  3733 => (x"86",x"c4",x"87",x"d8"),
  3734 => (x"fe",x"49",x"4c",x"73"),
  3735 => (x"70",x"87",x"f8",x"f0"),
  3736 => (x"87",x"cc",x"05",x"98"),
  3737 => (x"f0",x"fe",x"49",x"74"),
  3738 => (x"98",x"70",x"87",x"ed"),
  3739 => (x"87",x"f4",x"ff",x"02"),
  3740 => (x"e2",x"fe",x"49",x"c0"),
  3741 => (x"49",x"75",x"87",x"f0"),
  3742 => (x"87",x"fe",x"c9",x"fe"),
  3743 => (x"99",x"c2",x"49",x"70"),
  3744 => (x"c1",x"87",x"d4",x"05"),
  3745 => (x"eb",x"c6",x"fe",x"49"),
  3746 => (x"fe",x"49",x"75",x"87"),
  3747 => (x"70",x"87",x"eb",x"c9"),
  3748 => (x"02",x"99",x"c2",x"49"),
  3749 => (x"75",x"87",x"ec",x"ff"),
  3750 => (x"dd",x"c9",x"fe",x"49"),
  3751 => (x"02",x"98",x"70",x"87"),
  3752 => (x"c1",x"87",x"d2",x"c0"),
  3753 => (x"cb",x"c6",x"fe",x"49"),
  3754 => (x"fe",x"49",x"75",x"87"),
  3755 => (x"70",x"87",x"cb",x"c9"),
  3756 => (x"ee",x"ff",x"05",x"98"),
  3757 => (x"1e",x"e8",x"cf",x"87"),
  3758 => (x"49",x"d3",x"eb",x"c3"),
  3759 => (x"87",x"ee",x"ed",x"fe"),
  3760 => (x"c3",x"fc",x"86",x"c4"),
  3761 => (x"fb",x"e5",x"26",x"87"),
  3762 => (x"75",x"61",x"50",x"87"),
  3763 => (x"67",x"6e",x"69",x"73"),
  3764 => (x"55",x"00",x"2e",x"2e"),
  3765 => (x"75",x"61",x"70",x"6e"),
  3766 => (x"67",x"6e",x"69",x"73"),
  3767 => (x"00",x"2e",x"2e",x"2e"),
  3768 => (x"c8",x"d0",x"cb",x"cd"),
  3769 => (x"3e",x"3d",x"3c",x"3b"),
  3770 => (x"42",x"41",x"40",x"3f"),
  3771 => (x"00",x"d2",x"00",x"0e"),
  3772 => (x"00",x"9c",x"00",x"1c"),
  3773 => (x"08",x"9d",x"80",x"00"),
  3774 => (x"00",x"58",x"80",x"05"),
  3775 => (x"00",x"43",x"80",x"02"),
  3776 => (x"00",x"44",x"80",x"03"),
  3777 => (x"00",x"57",x"80",x"04"),
  3778 => (x"08",x"b8",x"80",x"01"),
  3779 => (x"00",x"00",x"00",x"04"),
  3780 => (x"00",x"00",x"00",x"11"),
  3781 => (x"00",x"00",x"00",x"1e"),
  3782 => (x"00",x"00",x"00",x"05"),
  3783 => (x"00",x"00",x"00",x"2c"),
  3784 => (x"00",x"00",x"00",x"1f"),
  3785 => (x"00",x"00",x"00",x"12"),
  3786 => (x"00",x"00",x"01",x"2a"),
  3787 => (x"00",x"00",x"00",x"06"),
  3788 => (x"00",x"00",x"00",x"13"),
  3789 => (x"00",x"00",x"00",x"20"),
  3790 => (x"00",x"00",x"00",x"07"),
  3791 => (x"00",x"00",x"00",x"2e"),
  3792 => (x"00",x"00",x"00",x"21"),
  3793 => (x"00",x"00",x"00",x"14"),
  3794 => (x"00",x"00",x"00",x"2d"),
  3795 => (x"00",x"47",x"00",x"08"),
  3796 => (x"00",x"00",x"00",x"15"),
  3797 => (x"00",x"00",x"00",x"22"),
  3798 => (x"00",x"48",x"00",x"09"),
  3799 => (x"00",x"00",x"00",x"30"),
  3800 => (x"00",x"00",x"00",x"23"),
  3801 => (x"00",x"4b",x"00",x"16"),
  3802 => (x"00",x"00",x"00",x"2f"),
  3803 => (x"00",x"49",x"00",x"0a"),
  3804 => (x"00",x"4c",x"00",x"17"),
  3805 => (x"00",x"4f",x"00",x"24"),
  3806 => (x"00",x"b5",x"00",x"0b"),
  3807 => (x"00",x"52",x"00",x"32"),
  3808 => (x"00",x"50",x"00",x"25"),
  3809 => (x"00",x"4d",x"00",x"18"),
  3810 => (x"00",x"00",x"00",x"31"),
  3811 => (x"00",x"00",x"00",x"0d"),
  3812 => (x"00",x"37",x"00",x"19"),
  3813 => (x"00",x"51",x"00",x"26"),
  3814 => (x"00",x"00",x"00",x"0c"),
  3815 => (x"00",x"53",x"00",x"34"),
  3816 => (x"00",x"4a",x"00",x"27"),
  3817 => (x"00",x"45",x"00",x"1a"),
  3818 => (x"00",x"00",x"00",x"33"),
  3819 => (x"00",x"cf",x"00",x"42"),
  3820 => (x"00",x"37",x"00",x"1b"),
  3821 => (x"00",x"00",x"00",x"28"),
  3822 => (x"00",x"c7",x"00",x"d3"),
  3823 => (x"00",x"00",x"02",x"36"),
  3824 => (x"00",x"2b",x"00",x"29"),
  3825 => (x"00",x"00",x"00",x"2b"),
  3826 => (x"00",x"4e",x"00",x"35"),
  3827 => (x"00",x"45",x"00",x"02"),
  3828 => (x"00",x"58",x"00",x"01"),
  3829 => (x"00",x"0f",x"04",x"1d"),
  3830 => (x"00",x"00",x"00",x"03"),
  3831 => (x"00",x"00",x"00",x"39"),
  3832 => (x"00",x"00",x"00",x"38"),
  3833 => (x"00",x"00",x"00",x"10"),
  3834 => (x"00",x"00",x"40",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

