///////////////   GLOBAL DEFINES   ////////////////
	
`define GUEST_TOP Next186_MiST	// substitute guest_top (lowercase) by guest's Mist top module name		

