library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"cccfc487",
    12 => x"86c0c64e",
    13 => x"49cccfc4",
    14 => x"48ecefc3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e6e7",
    19 => x"1e87fc98",
    20 => x"4a7186fc",
    21 => x"6949c0ff",
    22 => x"98c0c448",
    23 => x"026e7e70",
    24 => x"797287f5",
    25 => x"268efc48",
    26 => x"5b5e0e4f",
    27 => x"4b710e5c",
    28 => x"4a134cc0",
    29 => x"87cd029a",
    30 => x"d2ff4972",
    31 => x"1384c187",
    32 => x"f3059a4a",
    33 => x"26487487",
    34 => x"264b264c",
    35 => x"1e721e4f",
    36 => x"48121e73",
    37 => x"87ca0211",
    38 => x"98dfc34b",
    39 => x"0288739b",
    40 => x"4b2687f0",
    41 => x"4f264a26",
    42 => x"721e731e",
    43 => x"048bc11e",
    44 => x"481287ca",
    45 => x"87c40211",
    46 => x"87f10288",
    47 => x"4b264a26",
    48 => x"741e4f26",
    49 => x"721e731e",
    50 => x"048bc11e",
    51 => x"481287d0",
    52 => x"87ca0211",
    53 => x"98dfc34c",
    54 => x"0288749c",
    55 => x"4a2687eb",
    56 => x"4c264b26",
    57 => x"731e4f26",
    58 => x"a9738148",
    59 => x"1287c502",
    60 => x"87f60553",
    61 => x"c41e4f26",
    62 => x"48714a66",
    63 => x"fb055112",
    64 => x"1e4f2687",
    65 => x"73814873",
    66 => x"537205a9",
    67 => x"4f2687f9",
    68 => x"721e731e",
    69 => x"e7c0029a",
    70 => x"c148c087",
    71 => x"06a9724b",
    72 => x"827287d1",
    73 => x"7387c906",
    74 => x"01a97283",
    75 => x"87c387f4",
    76 => x"723ab2c1",
    77 => x"738903a9",
    78 => x"2ac10780",
    79 => x"87f3052b",
    80 => x"4f264b26",
    81 => x"c41e751e",
    82 => x"a1b7714d",
    83 => x"c1b9ff04",
    84 => x"07bdc381",
    85 => x"04a2b772",
    86 => x"82c1baff",
    87 => x"fe07bdc1",
    88 => x"2dc187ee",
    89 => x"c1b8ff04",
    90 => x"042d0780",
    91 => x"81c1b9ff",
    92 => x"264d2607",
    93 => x"48111e4f",
    94 => x"7808d4ff",
    95 => x"c14866c4",
    96 => x"58a6c888",
    97 => x"ed059870",
    98 => x"1e4f2687",
    99 => x"c348d4ff",
   100 => x"516878ff",
   101 => x"c14866c4",
   102 => x"58a6c888",
   103 => x"eb059870",
   104 => x"1e4f2687",
   105 => x"d4ff1e73",
   106 => x"7bffc34b",
   107 => x"ffc34a6b",
   108 => x"c8496b7b",
   109 => x"c3b17232",
   110 => x"4a6b7bff",
   111 => x"b27131c8",
   112 => x"6b7bffc3",
   113 => x"7232c849",
   114 => x"c44871b1",
   115 => x"264d2687",
   116 => x"264b264c",
   117 => x"5b5e0e4f",
   118 => x"710e5d5c",
   119 => x"4cd4ff4a",
   120 => x"ffc34972",
   121 => x"c37c7199",
   122 => x"05bfecef",
   123 => x"66d087c8",
   124 => x"d430c948",
   125 => x"66d058a6",
   126 => x"c329d849",
   127 => x"7c7199ff",
   128 => x"d04966d0",
   129 => x"99ffc329",
   130 => x"66d07c71",
   131 => x"c329c849",
   132 => x"7c7199ff",
   133 => x"c34966d0",
   134 => x"7c7199ff",
   135 => x"29d04972",
   136 => x"7199ffc3",
   137 => x"c94b6c7c",
   138 => x"c34dfff0",
   139 => x"d005abff",
   140 => x"7cffc387",
   141 => x"8dc14b6c",
   142 => x"c387c602",
   143 => x"f002abff",
   144 => x"fe487387",
   145 => x"c01e87c7",
   146 => x"48d4ff49",
   147 => x"c178ffc3",
   148 => x"b7c8c381",
   149 => x"87f104a9",
   150 => x"731e4f26",
   151 => x"c487e71e",
   152 => x"c04bdff8",
   153 => x"f0ffc01e",
   154 => x"fd49f7c1",
   155 => x"86c487e7",
   156 => x"c005a8c1",
   157 => x"d4ff87ea",
   158 => x"78ffc348",
   159 => x"c0c0c0c1",
   160 => x"c01ec0c0",
   161 => x"e9c1f0e1",
   162 => x"87c9fd49",
   163 => x"987086c4",
   164 => x"ff87ca05",
   165 => x"ffc348d4",
   166 => x"cb48c178",
   167 => x"87e6fe87",
   168 => x"fe058bc1",
   169 => x"48c087fd",
   170 => x"1e87e6fc",
   171 => x"d4ff1e73",
   172 => x"78ffc348",
   173 => x"1ec04bd3",
   174 => x"c1f0ffc0",
   175 => x"d4fc49c1",
   176 => x"7086c487",
   177 => x"87ca0598",
   178 => x"c348d4ff",
   179 => x"48c178ff",
   180 => x"f1fd87cb",
   181 => x"058bc187",
   182 => x"c087dbff",
   183 => x"87f1fb48",
   184 => x"5c5b5e0e",
   185 => x"4cd4ff0e",
   186 => x"c687dbfd",
   187 => x"e1c01eea",
   188 => x"49c8c1f0",
   189 => x"c487defb",
   190 => x"02a8c186",
   191 => x"eafe87c8",
   192 => x"c148c087",
   193 => x"dafa87e2",
   194 => x"cf497087",
   195 => x"c699ffff",
   196 => x"c802a9ea",
   197 => x"87d3fe87",
   198 => x"cbc148c0",
   199 => x"7cffc387",
   200 => x"fc4bf1c0",
   201 => x"987087f4",
   202 => x"87ebc002",
   203 => x"ffc01ec0",
   204 => x"49fac1f0",
   205 => x"c487defa",
   206 => x"05987086",
   207 => x"ffc387d9",
   208 => x"c3496c7c",
   209 => x"7c7c7cff",
   210 => x"99c0c17c",
   211 => x"c187c402",
   212 => x"c087d548",
   213 => x"c287d148",
   214 => x"87c405ab",
   215 => x"87c848c0",
   216 => x"fe058bc1",
   217 => x"48c087fd",
   218 => x"1e87e4f9",
   219 => x"efc31e73",
   220 => x"78c148ec",
   221 => x"d0ff4bc7",
   222 => x"fb78c248",
   223 => x"d0ff87c8",
   224 => x"c078c348",
   225 => x"d0e5c01e",
   226 => x"f949c0c1",
   227 => x"86c487c7",
   228 => x"c105a8c1",
   229 => x"abc24b87",
   230 => x"c087c505",
   231 => x"87f9c048",
   232 => x"ff058bc1",
   233 => x"f7fc87d0",
   234 => x"f0efc387",
   235 => x"05987058",
   236 => x"1ec187cd",
   237 => x"c1f0ffc0",
   238 => x"d8f849d0",
   239 => x"ff86c487",
   240 => x"ffc348d4",
   241 => x"87e0c478",
   242 => x"58f4efc3",
   243 => x"c248d0ff",
   244 => x"48d4ff78",
   245 => x"c178ffc3",
   246 => x"87f5f748",
   247 => x"5c5b5e0e",
   248 => x"4a710e5d",
   249 => x"ff4dffc3",
   250 => x"7c754cd4",
   251 => x"c448d0ff",
   252 => x"7c7578c3",
   253 => x"ffc01e72",
   254 => x"49d8c1f0",
   255 => x"c487d6f7",
   256 => x"02987086",
   257 => x"48c087c5",
   258 => x"7587f0c0",
   259 => x"7cfec37c",
   260 => x"d41ec0c8",
   261 => x"dcf54966",
   262 => x"7586c487",
   263 => x"757c757c",
   264 => x"e0dad87c",
   265 => x"6c7c754b",
   266 => x"c5059949",
   267 => x"058bc187",
   268 => x"7c7587f3",
   269 => x"c248d0ff",
   270 => x"f648c178",
   271 => x"ff1e87cf",
   272 => x"d0ff4ad4",
   273 => x"78d1c448",
   274 => x"c17affc3",
   275 => x"87f80589",
   276 => x"731e4f26",
   277 => x"c54b711e",
   278 => x"4adfcdee",
   279 => x"c348d4ff",
   280 => x"486878ff",
   281 => x"02a8fec3",
   282 => x"8ac187c5",
   283 => x"7287ed05",
   284 => x"87c5059a",
   285 => x"eac048c0",
   286 => x"029b7387",
   287 => x"66c887cc",
   288 => x"f449731e",
   289 => x"86c487c5",
   290 => x"66c887c6",
   291 => x"87eefe49",
   292 => x"c348d4ff",
   293 => x"737878ff",
   294 => x"87c5059b",
   295 => x"d048d0ff",
   296 => x"f448c178",
   297 => x"731e87eb",
   298 => x"c04a711e",
   299 => x"48d4ff4b",
   300 => x"ff78ffc3",
   301 => x"c3c448d0",
   302 => x"48d4ff78",
   303 => x"7278ffc3",
   304 => x"f0ffc01e",
   305 => x"f449d1c1",
   306 => x"86c487cb",
   307 => x"cd059870",
   308 => x"1ec0c887",
   309 => x"fd4966cc",
   310 => x"86c487f8",
   311 => x"d0ff4b70",
   312 => x"7378c248",
   313 => x"87e9f348",
   314 => x"5c5b5e0e",
   315 => x"1ec00e5d",
   316 => x"c1f0ffc0",
   317 => x"dcf349c9",
   318 => x"c31ed287",
   319 => x"fd49f4ef",
   320 => x"86c887d0",
   321 => x"84c14cc0",
   322 => x"04acb7d2",
   323 => x"efc387f8",
   324 => x"49bf97f4",
   325 => x"c199c0c3",
   326 => x"c005a9c0",
   327 => x"efc387e7",
   328 => x"49bf97fb",
   329 => x"efc331d0",
   330 => x"4abf97fc",
   331 => x"b17232c8",
   332 => x"97fdefc3",
   333 => x"71b14abf",
   334 => x"ffffcf4c",
   335 => x"84c19cff",
   336 => x"e7c134ca",
   337 => x"fdefc387",
   338 => x"c149bf97",
   339 => x"c399c631",
   340 => x"bf97feef",
   341 => x"2ab7c74a",
   342 => x"efc3b172",
   343 => x"4abf97f9",
   344 => x"c39dcf4d",
   345 => x"bf97faef",
   346 => x"ca9ac34a",
   347 => x"fbefc332",
   348 => x"c24bbf97",
   349 => x"c3b27333",
   350 => x"bf97fcef",
   351 => x"9bc0c34b",
   352 => x"732bb7c6",
   353 => x"c181c2b2",
   354 => x"70307148",
   355 => x"7548c149",
   356 => x"724d7030",
   357 => x"7184c14c",
   358 => x"b7c0c894",
   359 => x"87cc06ad",
   360 => x"2db734c1",
   361 => x"adb7c0c8",
   362 => x"87f4ff01",
   363 => x"dcf04874",
   364 => x"5b5e0e87",
   365 => x"f80e5d5c",
   366 => x"daf8c386",
   367 => x"c378c048",
   368 => x"c01ed2f0",
   369 => x"87defb49",
   370 => x"987086c4",
   371 => x"c087c505",
   372 => x"87cec948",
   373 => x"7ec14dc0",
   374 => x"bff0fbc0",
   375 => x"c8f1c349",
   376 => x"4bc8714a",
   377 => x"7087c1eb",
   378 => x"87c20598",
   379 => x"fbc07ec0",
   380 => x"c349bfec",
   381 => x"714ae4f1",
   382 => x"ebea4bc8",
   383 => x"05987087",
   384 => x"7ec087c2",
   385 => x"fdc0026e",
   386 => x"d8f7c387",
   387 => x"f8c34dbf",
   388 => x"7ebf9fd0",
   389 => x"ead6c548",
   390 => x"87c705a8",
   391 => x"bfd8f7c3",
   392 => x"6e87ce4d",
   393 => x"d5e9ca48",
   394 => x"87c502a8",
   395 => x"f1c748c0",
   396 => x"d2f0c387",
   397 => x"f949751e",
   398 => x"86c487ec",
   399 => x"c5059870",
   400 => x"c748c087",
   401 => x"fbc087dc",
   402 => x"c349bfec",
   403 => x"714ae4f1",
   404 => x"d3e94bc8",
   405 => x"05987087",
   406 => x"f8c387c8",
   407 => x"78c148da",
   408 => x"fbc087da",
   409 => x"c349bff0",
   410 => x"714ac8f1",
   411 => x"f7e84bc8",
   412 => x"02987087",
   413 => x"c087c5c0",
   414 => x"87e6c648",
   415 => x"97d0f8c3",
   416 => x"d5c149bf",
   417 => x"cdc005a9",
   418 => x"d1f8c387",
   419 => x"c249bf97",
   420 => x"c002a9ea",
   421 => x"48c087c5",
   422 => x"c387c7c6",
   423 => x"bf97d2f0",
   424 => x"e9c3487e",
   425 => x"cec002a8",
   426 => x"c3486e87",
   427 => x"c002a8eb",
   428 => x"48c087c5",
   429 => x"c387ebc5",
   430 => x"bf97ddf0",
   431 => x"c0059949",
   432 => x"f0c387cc",
   433 => x"49bf97de",
   434 => x"c002a9c2",
   435 => x"48c087c5",
   436 => x"c387cfc5",
   437 => x"bf97dff0",
   438 => x"d6f8c348",
   439 => x"484c7058",
   440 => x"f8c388c1",
   441 => x"f0c358da",
   442 => x"49bf97e0",
   443 => x"f0c38175",
   444 => x"4abf97e1",
   445 => x"a17232c8",
   446 => x"e7fcc37e",
   447 => x"c3786e48",
   448 => x"bf97e2f0",
   449 => x"58a6c848",
   450 => x"bfdaf8c3",
   451 => x"87d4c202",
   452 => x"bfecfbc0",
   453 => x"e4f1c349",
   454 => x"4bc8714a",
   455 => x"7087c9e6",
   456 => x"c5c00298",
   457 => x"c348c087",
   458 => x"f8c387f8",
   459 => x"c34cbfd2",
   460 => x"c35cfbfc",
   461 => x"bf97f7f0",
   462 => x"c331c849",
   463 => x"bf97f6f0",
   464 => x"c349a14a",
   465 => x"bf97f8f0",
   466 => x"7232d04a",
   467 => x"f0c349a1",
   468 => x"4abf97f9",
   469 => x"a17232d8",
   470 => x"9166c449",
   471 => x"bfe7fcc3",
   472 => x"effcc381",
   473 => x"fff0c359",
   474 => x"c84abf97",
   475 => x"fef0c332",
   476 => x"a24bbf97",
   477 => x"c0f1c34a",
   478 => x"d04bbf97",
   479 => x"4aa27333",
   480 => x"97c1f1c3",
   481 => x"9bcf4bbf",
   482 => x"a27333d8",
   483 => x"f3fcc34a",
   484 => x"effcc35a",
   485 => x"8ac24abf",
   486 => x"fcc39274",
   487 => x"a17248f3",
   488 => x"87cac178",
   489 => x"97e4f0c3",
   490 => x"31c849bf",
   491 => x"97e3f0c3",
   492 => x"49a14abf",
   493 => x"59e2f8c3",
   494 => x"bfdef8c3",
   495 => x"c731c549",
   496 => x"29c981ff",
   497 => x"59fbfcc3",
   498 => x"97e9f0c3",
   499 => x"32c84abf",
   500 => x"97e8f0c3",
   501 => x"4aa24bbf",
   502 => x"6e9266c4",
   503 => x"f7fcc382",
   504 => x"effcc35a",
   505 => x"c378c048",
   506 => x"7248ebfc",
   507 => x"fcc378a1",
   508 => x"fcc348fb",
   509 => x"c378bfef",
   510 => x"c348fffc",
   511 => x"78bff3fc",
   512 => x"bfdaf8c3",
   513 => x"87c9c002",
   514 => x"30c44874",
   515 => x"c9c07e70",
   516 => x"f7fcc387",
   517 => x"30c448bf",
   518 => x"f8c37e70",
   519 => x"786e48de",
   520 => x"8ef848c1",
   521 => x"4c264d26",
   522 => x"4f264b26",
   523 => x"5c5b5e0e",
   524 => x"4a710e5d",
   525 => x"bfdaf8c3",
   526 => x"7287cb02",
   527 => x"722bc74b",
   528 => x"9cffc14c",
   529 => x"4b7287c9",
   530 => x"4c722bc8",
   531 => x"c39cffc3",
   532 => x"83bfe7fc",
   533 => x"bfe8fbc0",
   534 => x"87d902ab",
   535 => x"5becfbc0",
   536 => x"1ed2f0c3",
   537 => x"fdf04973",
   538 => x"7086c487",
   539 => x"87c50598",
   540 => x"e6c048c0",
   541 => x"daf8c387",
   542 => x"87d202bf",
   543 => x"91c44974",
   544 => x"81d2f0c3",
   545 => x"ffcf4d69",
   546 => x"9dffffff",
   547 => x"497487cb",
   548 => x"f0c391c2",
   549 => x"699f81d2",
   550 => x"fe48754d",
   551 => x"5e0e87c6",
   552 => x"0e5d5c5b",
   553 => x"c04d711e",
   554 => x"d149c11e",
   555 => x"86c487e2",
   556 => x"029c4c70",
   557 => x"c387c2c1",
   558 => x"754ae2f8",
   559 => x"ccdfff49",
   560 => x"02987087",
   561 => x"7487f2c0",
   562 => x"cb49754a",
   563 => x"f1dfff4b",
   564 => x"02987087",
   565 => x"c087e2c0",
   566 => x"029c741e",
   567 => x"a6c487c7",
   568 => x"c578c048",
   569 => x"48a6c487",
   570 => x"66c478c1",
   571 => x"87e0d049",
   572 => x"4c7086c4",
   573 => x"fefe059c",
   574 => x"26487487",
   575 => x"0e87e5fc",
   576 => x"5d5c5b5e",
   577 => x"7186f80e",
   578 => x"c5059b4b",
   579 => x"c248c087",
   580 => x"a3c887d4",
   581 => x"d87dc04d",
   582 => x"87c70266",
   583 => x"bf9766d8",
   584 => x"c087c505",
   585 => x"87fec148",
   586 => x"fd4966d8",
   587 => x"7e7087f0",
   588 => x"efc1026e",
   589 => x"dc496e87",
   590 => x"6e7d6981",
   591 => x"c481da49",
   592 => x"699f4ca3",
   593 => x"daf8c37c",
   594 => x"87d002bf",
   595 => x"81d4496e",
   596 => x"4a49699f",
   597 => x"9affffc0",
   598 => x"87c232d0",
   599 => x"49724ac0",
   600 => x"70806c48",
   601 => x"cc7bc07c",
   602 => x"796c49a3",
   603 => x"c049a3d0",
   604 => x"48a6c479",
   605 => x"a3d478c0",
   606 => x"4966c44a",
   607 => x"a17291c8",
   608 => x"6c41c049",
   609 => x"4866c479",
   610 => x"a6c880c1",
   611 => x"a8b7d058",
   612 => x"87e2ff04",
   613 => x"2ac94a6d",
   614 => x"d4c22ac7",
   615 => x"797249a3",
   616 => x"87c2486e",
   617 => x"8ef848c0",
   618 => x"0e87f9f9",
   619 => x"5d5c5b5e",
   620 => x"c04c710e",
   621 => x"ff48e8fb",
   622 => x"029c7478",
   623 => x"c887cac1",
   624 => x"026949a4",
   625 => x"d087c2c1",
   626 => x"496c4a66",
   627 => x"5aa6d482",
   628 => x"b94d66d0",
   629 => x"bfd6f8c3",
   630 => x"72baff4a",
   631 => x"02997199",
   632 => x"c487e4c0",
   633 => x"496b4ba4",
   634 => x"7087c1f9",
   635 => x"d2f8c37b",
   636 => x"816c49bf",
   637 => x"b9757c71",
   638 => x"bfd6f8c3",
   639 => x"72baff4a",
   640 => x"05997199",
   641 => x"7587dcff",
   642 => x"87d8f87c",
   643 => x"711e731e",
   644 => x"c7029b4b",
   645 => x"49a3c887",
   646 => x"87c50569",
   647 => x"ebc048c0",
   648 => x"ebfcc387",
   649 => x"a3c44abf",
   650 => x"c2496949",
   651 => x"d2f8c389",
   652 => x"a27191bf",
   653 => x"d6f8c34a",
   654 => x"996b49bf",
   655 => x"c84aa271",
   656 => x"49721e66",
   657 => x"c487dfe9",
   658 => x"48497086",
   659 => x"1e87d9f7",
   660 => x"4b711e73",
   661 => x"87c7029b",
   662 => x"6949a3c8",
   663 => x"c087c505",
   664 => x"87ebc048",
   665 => x"bfebfcc3",
   666 => x"49a3c44a",
   667 => x"89c24969",
   668 => x"bfd2f8c3",
   669 => x"4aa27191",
   670 => x"bfd6f8c3",
   671 => x"71996b49",
   672 => x"66c84aa2",
   673 => x"e549721e",
   674 => x"86c487d2",
   675 => x"f6484970",
   676 => x"5e0e87d6",
   677 => x"0e5d5c5b",
   678 => x"4b7186f8",
   679 => x"ff48a6c4",
   680 => x"49a3c878",
   681 => x"4cc04d69",
   682 => x"744aa3d4",
   683 => x"7291c849",
   684 => x"496949a1",
   685 => x"714866d8",
   686 => x"d87e7088",
   687 => x"ca01a966",
   688 => x"06ad6e87",
   689 => x"a6c887c5",
   690 => x"c14d6e5c",
   691 => x"acb7d084",
   692 => x"87d4ff04",
   693 => x"f84866c4",
   694 => x"87c8f58e",
   695 => x"5c5b5e0e",
   696 => x"86ec0e5d",
   697 => x"c859a6c8",
   698 => x"ffc148a6",
   699 => x"ffffffff",
   700 => x"ff80c478",
   701 => x"c04dc078",
   702 => x"4b66c44c",
   703 => x"497483d4",
   704 => x"a17391c8",
   705 => x"c84a7549",
   706 => x"7ea27392",
   707 => x"bf6e4969",
   708 => x"59a6d489",
   709 => x"c605ad74",
   710 => x"48a6d087",
   711 => x"d078bf6e",
   712 => x"b7c04866",
   713 => x"87cf04a8",
   714 => x"c84966d0",
   715 => x"c603a966",
   716 => x"5ca6d087",
   717 => x"c159a6cc",
   718 => x"acb7d084",
   719 => x"87f9fe04",
   720 => x"b7d085c1",
   721 => x"eefe04ad",
   722 => x"4866cc87",
   723 => x"d3f38eec",
   724 => x"5b5e0e87",
   725 => x"4b710e5c",
   726 => x"a3c84cc0",
   727 => x"c4496949",
   728 => x"914a7429",
   729 => x"49731e71",
   730 => x"86c487d4",
   731 => x"b7d084c1",
   732 => x"87e604ac",
   733 => x"49731ec0",
   734 => x"f22687c4",
   735 => x"5e0e87e8",
   736 => x"0e5d5c5b",
   737 => x"4b7186f0",
   738 => x"4c66e0c0",
   739 => x"9b732cc9",
   740 => x"87e1c302",
   741 => x"6949a3c8",
   742 => x"87d9c302",
   743 => x"c049a3d0",
   744 => x"6b7966e0",
   745 => x"c302ac7e",
   746 => x"f8c387cb",
   747 => x"ff49bfd6",
   748 => x"744a71b9",
   749 => x"6e48719a",
   750 => x"58a6cc98",
   751 => x"c44da3c4",
   752 => x"786d48a6",
   753 => x"05aa66c8",
   754 => x"7b7487c5",
   755 => x"7287d1c2",
   756 => x"fa49731e",
   757 => x"86c487fc",
   758 => x"c0487e70",
   759 => x"d004a8b7",
   760 => x"4aa3d487",
   761 => x"91c8496e",
   762 => x"2149a172",
   763 => x"c77d697b",
   764 => x"cc7bc087",
   765 => x"7d6949a3",
   766 => x"731e66c8",
   767 => x"87d2fa49",
   768 => x"7e7086c4",
   769 => x"49a3d4c2",
   770 => x"6948a6cc",
   771 => x"4866c878",
   772 => x"06a866cc",
   773 => x"486e87c9",
   774 => x"04a8b7c0",
   775 => x"6e87e0c0",
   776 => x"a8b7c048",
   777 => x"87ecc004",
   778 => x"6e4aa3d4",
   779 => x"7291c849",
   780 => x"66c849a1",
   781 => x"70886948",
   782 => x"a966cc49",
   783 => x"7387d506",
   784 => x"87d8fa49",
   785 => x"a3d44970",
   786 => x"7291c84a",
   787 => x"66c849a1",
   788 => x"7966c441",
   789 => x"49748c6b",
   790 => x"f549731e",
   791 => x"86c487cd",
   792 => x"4966e0c0",
   793 => x"0299ffc7",
   794 => x"f0c387cb",
   795 => x"49731ed2",
   796 => x"c487d9f6",
   797 => x"ee8ef086",
   798 => x"731e87ea",
   799 => x"9b4b711e",
   800 => x"87e4c002",
   801 => x"5bfffcc3",
   802 => x"8ac24a73",
   803 => x"bfd2f8c3",
   804 => x"fcc39249",
   805 => x"7248bfeb",
   806 => x"c3fdc380",
   807 => x"c4487158",
   808 => x"e2f8c330",
   809 => x"87edc058",
   810 => x"48fbfcc3",
   811 => x"bfeffcc3",
   812 => x"fffcc378",
   813 => x"f3fcc348",
   814 => x"f8c378bf",
   815 => x"c902bfda",
   816 => x"d2f8c387",
   817 => x"31c449bf",
   818 => x"fcc387c7",
   819 => x"c449bff7",
   820 => x"e2f8c331",
   821 => x"87d0ed59",
   822 => x"5c5b5e0e",
   823 => x"c04a710e",
   824 => x"029a724b",
   825 => x"da87e1c0",
   826 => x"699f49a2",
   827 => x"daf8c34b",
   828 => x"87cf02bf",
   829 => x"9f49a2d4",
   830 => x"c04c4969",
   831 => x"d09cffff",
   832 => x"c087c234",
   833 => x"b349744c",
   834 => x"edfd4973",
   835 => x"87d6ec87",
   836 => x"5c5b5e0e",
   837 => x"86f40e5d",
   838 => x"7ec04a71",
   839 => x"d8029a72",
   840 => x"cef0c387",
   841 => x"c378c048",
   842 => x"c348c6f0",
   843 => x"78bffffc",
   844 => x"48caf0c3",
   845 => x"bffbfcc3",
   846 => x"eff8c378",
   847 => x"c350c048",
   848 => x"49bfdef8",
   849 => x"bfcef0c3",
   850 => x"03aa714a",
   851 => x"7287c0c4",
   852 => x"0599cf49",
   853 => x"c387e1c0",
   854 => x"c31ed2f0",
   855 => x"49bfc6f0",
   856 => x"48c6f0c3",
   857 => x"7178a1c1",
   858 => x"87fadcff",
   859 => x"fbc086c4",
   860 => x"f0c348e4",
   861 => x"87cc78d2",
   862 => x"bfe4fbc0",
   863 => x"80e0c048",
   864 => x"58e8fbc0",
   865 => x"bfcef0c3",
   866 => x"c380c148",
   867 => x"2758d2f0",
   868 => x"00000ee4",
   869 => x"4dbf97bf",
   870 => x"e2c2029d",
   871 => x"ade5c387",
   872 => x"87dbc202",
   873 => x"bfe4fbc0",
   874 => x"49a3cb4b",
   875 => x"accf4c11",
   876 => x"87d2c105",
   877 => x"99df4975",
   878 => x"91cd89c1",
   879 => x"81e2f8c3",
   880 => x"124aa3c1",
   881 => x"4aa3c351",
   882 => x"a3c55112",
   883 => x"c751124a",
   884 => x"51124aa3",
   885 => x"124aa3c9",
   886 => x"4aa3ce51",
   887 => x"a3d05112",
   888 => x"d251124a",
   889 => x"51124aa3",
   890 => x"124aa3d4",
   891 => x"4aa3d651",
   892 => x"a3d85112",
   893 => x"dc51124a",
   894 => x"51124aa3",
   895 => x"124aa3de",
   896 => x"c07ec151",
   897 => x"497487f9",
   898 => x"c00599c8",
   899 => x"497487ea",
   900 => x"d00599d0",
   901 => x"0266dc87",
   902 => x"7387cac0",
   903 => x"0f66dc49",
   904 => x"d3029870",
   905 => x"c0056e87",
   906 => x"f8c387c6",
   907 => x"50c048e2",
   908 => x"bfe4fbc0",
   909 => x"87e7c248",
   910 => x"48eff8c3",
   911 => x"c37e50c0",
   912 => x"49bfdef8",
   913 => x"bfcef0c3",
   914 => x"04aa714a",
   915 => x"c387c0fc",
   916 => x"05bffffc",
   917 => x"c387c8c0",
   918 => x"02bfdaf8",
   919 => x"c087fec1",
   920 => x"ff48e8fb",
   921 => x"caf0c378",
   922 => x"ffe649bf",
   923 => x"c3497087",
   924 => x"c459cef0",
   925 => x"f0c348a6",
   926 => x"c378bfca",
   927 => x"02bfdaf8",
   928 => x"c487d8c0",
   929 => x"ffcf4966",
   930 => x"99f8ffff",
   931 => x"c5c002a9",
   932 => x"c04dc087",
   933 => x"4dc187e1",
   934 => x"c487dcc0",
   935 => x"ffcf4966",
   936 => x"02a999f8",
   937 => x"c887c8c0",
   938 => x"78c048a6",
   939 => x"c887c5c0",
   940 => x"78c148a6",
   941 => x"754d66c8",
   942 => x"e0c0059d",
   943 => x"4966c487",
   944 => x"f8c389c2",
   945 => x"914abfd2",
   946 => x"bfebfcc3",
   947 => x"c6f0c34a",
   948 => x"78a17248",
   949 => x"48cef0c3",
   950 => x"e2f978c0",
   951 => x"f448c087",
   952 => x"87c0e58e",
   953 => x"00000000",
   954 => x"ffffffff",
   955 => x"00000ef4",
   956 => x"00000efd",
   957 => x"33544146",
   958 => x"20202032",
   959 => x"54414600",
   960 => x"20203631",
   961 => x"ff1e0020",
   962 => x"ffc348d4",
   963 => x"26486878",
   964 => x"d4ff1e4f",
   965 => x"78ffc348",
   966 => x"c848d0ff",
   967 => x"d4ff78e1",
   968 => x"c378d448",
   969 => x"ff48c3fd",
   970 => x"2650bfd4",
   971 => x"d0ff1e4f",
   972 => x"78e0c048",
   973 => x"ff1e4f26",
   974 => x"497087cc",
   975 => x"87c60299",
   976 => x"05a9fbc0",
   977 => x"487187f1",
   978 => x"5e0e4f26",
   979 => x"710e5c5b",
   980 => x"fe4cc04b",
   981 => x"497087f0",
   982 => x"f9c00299",
   983 => x"a9ecc087",
   984 => x"87f2c002",
   985 => x"02a9fbc0",
   986 => x"cc87ebc0",
   987 => x"03acb766",
   988 => x"66d087c7",
   989 => x"7187c202",
   990 => x"02997153",
   991 => x"84c187c2",
   992 => x"7087c3fe",
   993 => x"cd029949",
   994 => x"a9ecc087",
   995 => x"c087c702",
   996 => x"ff05a9fb",
   997 => x"66d087d5",
   998 => x"c087c302",
   999 => x"ecc07b97",
  1000 => x"87c405a9",
  1001 => x"87c54a74",
  1002 => x"0ac04a74",
  1003 => x"c248728a",
  1004 => x"264d2687",
  1005 => x"264b264c",
  1006 => x"c9fd1e4f",
  1007 => x"c0497087",
  1008 => x"04a9b7f0",
  1009 => x"f9c087ca",
  1010 => x"c301a9b7",
  1011 => x"89f0c087",
  1012 => x"a9b7c1c1",
  1013 => x"c187ca04",
  1014 => x"01a9b7da",
  1015 => x"f7c087c3",
  1016 => x"26487189",
  1017 => x"5b5e0e4f",
  1018 => x"4c710e5c",
  1019 => x"c187e2fc",
  1020 => x"1e66d01e",
  1021 => x"d1fd4974",
  1022 => x"7086c887",
  1023 => x"87edfc4b",
  1024 => x"03abb7c0",
  1025 => x"8b0b87c2",
  1026 => x"abb766cc",
  1027 => x"7487cf03",
  1028 => x"83c149a3",
  1029 => x"cc51e0c0",
  1030 => x"04abb766",
  1031 => x"a37487f1",
  1032 => x"fe51c049",
  1033 => x"5e0e87cd",
  1034 => x"710e5c5b",
  1035 => x"4cd4ff4a",
  1036 => x"eac04972",
  1037 => x"9b4b7087",
  1038 => x"c187c202",
  1039 => x"48d0ff8b",
  1040 => x"c178c5c8",
  1041 => x"49737cd5",
  1042 => x"cfc331c6",
  1043 => x"4abf97da",
  1044 => x"70b07148",
  1045 => x"48d0ff7c",
  1046 => x"487378c4",
  1047 => x"0e87d4fd",
  1048 => x"5d5c5b5e",
  1049 => x"7186f80e",
  1050 => x"fa7ec04c",
  1051 => x"4bc087e3",
  1052 => x"97ccc4c1",
  1053 => x"a9c049bf",
  1054 => x"fa87cf04",
  1055 => x"83c187f8",
  1056 => x"97ccc4c1",
  1057 => x"06ab49bf",
  1058 => x"c4c187f1",
  1059 => x"02bf97cc",
  1060 => x"f1f987cf",
  1061 => x"99497087",
  1062 => x"c087c602",
  1063 => x"f105a9ec",
  1064 => x"f94bc087",
  1065 => x"4d7087e0",
  1066 => x"c887dbf9",
  1067 => x"d5f958a6",
  1068 => x"c14a7087",
  1069 => x"49a4c883",
  1070 => x"ad496997",
  1071 => x"c087c702",
  1072 => x"c005adff",
  1073 => x"a4c987e7",
  1074 => x"49699749",
  1075 => x"02a966c4",
  1076 => x"c04887c7",
  1077 => x"d405a8ff",
  1078 => x"49a4ca87",
  1079 => x"aa496997",
  1080 => x"c087c602",
  1081 => x"c405aaff",
  1082 => x"d07ec187",
  1083 => x"adecc087",
  1084 => x"c087c602",
  1085 => x"c405adfb",
  1086 => x"c14bc087",
  1087 => x"fe026e7e",
  1088 => x"e8f887e1",
  1089 => x"f8487387",
  1090 => x"87e5fa8e",
  1091 => x"5b5e0e00",
  1092 => x"1e0e5d5c",
  1093 => x"4cc04b71",
  1094 => x"c004ab4d",
  1095 => x"c1c187e8",
  1096 => x"9d751edf",
  1097 => x"c087c402",
  1098 => x"c187c24a",
  1099 => x"ef49724a",
  1100 => x"86c487de",
  1101 => x"84c17e70",
  1102 => x"87c2056e",
  1103 => x"85c14c73",
  1104 => x"ff06ac73",
  1105 => x"486e87d8",
  1106 => x"264d2626",
  1107 => x"264b264c",
  1108 => x"5b5e0e4f",
  1109 => x"1e0e5d5c",
  1110 => x"de494c71",
  1111 => x"ddfdc391",
  1112 => x"9785714d",
  1113 => x"ddc1026d",
  1114 => x"c8fdc387",
  1115 => x"82744abf",
  1116 => x"d8fe4972",
  1117 => x"6e7e7087",
  1118 => x"87f3c002",
  1119 => x"4bd0fdc3",
  1120 => x"49cb4a6e",
  1121 => x"87defdfe",
  1122 => x"93cb4b74",
  1123 => x"83d7e9c1",
  1124 => x"c7c183c4",
  1125 => x"49747bca",
  1126 => x"87e5c4c1",
  1127 => x"fdc37b75",
  1128 => x"49bf97dc",
  1129 => x"d0fdc31e",
  1130 => x"c0dac249",
  1131 => x"7486c487",
  1132 => x"ccc4c149",
  1133 => x"c149c087",
  1134 => x"c387ebc5",
  1135 => x"c048c4fd",
  1136 => x"dd49c178",
  1137 => x"fd2687d1",
  1138 => x"6f4c87ff",
  1139 => x"6e696461",
  1140 => x"2e2e2e67",
  1141 => x"5b5e0e00",
  1142 => x"4b710e5c",
  1143 => x"c8fdc34a",
  1144 => x"497282bf",
  1145 => x"7087e6fc",
  1146 => x"c4029c4c",
  1147 => x"e7eb4987",
  1148 => x"c8fdc387",
  1149 => x"c178c048",
  1150 => x"87dbdc49",
  1151 => x"0e87ccfd",
  1152 => x"5d5c5b5e",
  1153 => x"c386f40e",
  1154 => x"c04dd2f0",
  1155 => x"48a6c44c",
  1156 => x"fdc378c0",
  1157 => x"c049bfc8",
  1158 => x"c1c106a9",
  1159 => x"d2f0c387",
  1160 => x"c0029848",
  1161 => x"c1c187f8",
  1162 => x"66c81edf",
  1163 => x"c487c702",
  1164 => x"78c048a6",
  1165 => x"a6c487c5",
  1166 => x"c478c148",
  1167 => x"cfeb4966",
  1168 => x"7086c487",
  1169 => x"c484c14d",
  1170 => x"80c14866",
  1171 => x"c358a6c8",
  1172 => x"49bfc8fd",
  1173 => x"87c603ac",
  1174 => x"ff059d75",
  1175 => x"4cc087c8",
  1176 => x"c3029d75",
  1177 => x"c1c187e0",
  1178 => x"66c81edf",
  1179 => x"cc87c702",
  1180 => x"78c048a6",
  1181 => x"a6cc87c5",
  1182 => x"cc78c148",
  1183 => x"cfea4966",
  1184 => x"7086c487",
  1185 => x"c2026e7e",
  1186 => x"496e87e9",
  1187 => x"699781cb",
  1188 => x"0299d049",
  1189 => x"c187d6c1",
  1190 => x"744ad5c7",
  1191 => x"c191cb49",
  1192 => x"7281d7e9",
  1193 => x"c381c879",
  1194 => x"497451ff",
  1195 => x"fdc391de",
  1196 => x"85714ddd",
  1197 => x"7d97c1c2",
  1198 => x"c049a5c1",
  1199 => x"f8c351e0",
  1200 => x"02bf97e2",
  1201 => x"84c187d2",
  1202 => x"c34ba5c2",
  1203 => x"db4ae2f8",
  1204 => x"d1f8fe49",
  1205 => x"87dbc187",
  1206 => x"c049a5cd",
  1207 => x"c284c151",
  1208 => x"4a6e4ba5",
  1209 => x"f7fe49cb",
  1210 => x"c6c187fc",
  1211 => x"d1c5c187",
  1212 => x"cb49744a",
  1213 => x"d7e9c191",
  1214 => x"c3797281",
  1215 => x"bf97e2f8",
  1216 => x"7487d802",
  1217 => x"c191de49",
  1218 => x"ddfdc384",
  1219 => x"c383714b",
  1220 => x"dd4ae2f8",
  1221 => x"cdf7fe49",
  1222 => x"7487d887",
  1223 => x"c393de4b",
  1224 => x"cb83ddfd",
  1225 => x"51c049a3",
  1226 => x"6e7384c1",
  1227 => x"fe49cb4a",
  1228 => x"c487f3f6",
  1229 => x"80c14866",
  1230 => x"c758a6c8",
  1231 => x"c5c003ac",
  1232 => x"fc056e87",
  1233 => x"487487e0",
  1234 => x"fcf78ef4",
  1235 => x"1e731e87",
  1236 => x"cb494b71",
  1237 => x"d7e9c191",
  1238 => x"4aa1c881",
  1239 => x"48dacfc3",
  1240 => x"a1c95012",
  1241 => x"ccc4c14a",
  1242 => x"ca501248",
  1243 => x"dcfdc381",
  1244 => x"c3501148",
  1245 => x"bf97dcfd",
  1246 => x"49c01e49",
  1247 => x"87edd2c2",
  1248 => x"48c4fdc3",
  1249 => x"49c178de",
  1250 => x"2687ccd6",
  1251 => x"1e87fef6",
  1252 => x"cb494a71",
  1253 => x"d7e9c191",
  1254 => x"1181c881",
  1255 => x"c8fdc348",
  1256 => x"c8fdc358",
  1257 => x"c178c048",
  1258 => x"87ebd549",
  1259 => x"c01e4f26",
  1260 => x"f1fdc049",
  1261 => x"1e4f2687",
  1262 => x"d2029971",
  1263 => x"eceac187",
  1264 => x"f750c048",
  1265 => x"cfcec180",
  1266 => x"d0e9c140",
  1267 => x"c187ce78",
  1268 => x"c148e8ea",
  1269 => x"fc78c9e9",
  1270 => x"eecec180",
  1271 => x"0e4f2678",
  1272 => x"0e5c5b5e",
  1273 => x"cb4a4c71",
  1274 => x"d7e9c192",
  1275 => x"49a2c882",
  1276 => x"974ba2c9",
  1277 => x"971e4b6b",
  1278 => x"ca1e4969",
  1279 => x"c0491282",
  1280 => x"c087ece8",
  1281 => x"87cfd449",
  1282 => x"fac04974",
  1283 => x"8ef887f3",
  1284 => x"1e87f8f4",
  1285 => x"4b711e73",
  1286 => x"87c3ff49",
  1287 => x"fefe4973",
  1288 => x"c049c087",
  1289 => x"f487fffb",
  1290 => x"731e87e3",
  1291 => x"c64b711e",
  1292 => x"db024aa3",
  1293 => x"028ac187",
  1294 => x"028a87d6",
  1295 => x"8a87dac1",
  1296 => x"87fcc002",
  1297 => x"e1c0028a",
  1298 => x"cb028a87",
  1299 => x"87dbc187",
  1300 => x"fafc49c7",
  1301 => x"87dec187",
  1302 => x"bfc8fdc3",
  1303 => x"87cbc102",
  1304 => x"c388c148",
  1305 => x"c158ccfd",
  1306 => x"fdc387c1",
  1307 => x"c002bfcc",
  1308 => x"fdc387f9",
  1309 => x"c148bfc8",
  1310 => x"ccfdc380",
  1311 => x"87ebc058",
  1312 => x"bfc8fdc3",
  1313 => x"c389c649",
  1314 => x"c059ccfd",
  1315 => x"da03a9b7",
  1316 => x"c8fdc387",
  1317 => x"d278c048",
  1318 => x"ccfdc387",
  1319 => x"87cb02bf",
  1320 => x"bfc8fdc3",
  1321 => x"c380c648",
  1322 => x"c058ccfd",
  1323 => x"87e7d149",
  1324 => x"f8c04973",
  1325 => x"d4f287cb",
  1326 => x"5b5e0e87",
  1327 => x"4c710e5c",
  1328 => x"741e66cc",
  1329 => x"c193cb4b",
  1330 => x"c483d7e9",
  1331 => x"496a4aa3",
  1332 => x"87e2f0fe",
  1333 => x"7bcdcdc1",
  1334 => x"d449a3c8",
  1335 => x"a3c95166",
  1336 => x"5166d849",
  1337 => x"dc49a3ca",
  1338 => x"f1265166",
  1339 => x"5e0e87dd",
  1340 => x"0e5d5c5b",
  1341 => x"d886d0ff",
  1342 => x"a6c459a6",
  1343 => x"c478c048",
  1344 => x"66c4c180",
  1345 => x"c180c478",
  1346 => x"c180c478",
  1347 => x"ccfdc378",
  1348 => x"c378c148",
  1349 => x"48bfc4fd",
  1350 => x"cb05a8de",
  1351 => x"87dff387",
  1352 => x"a6c84970",
  1353 => x"87f8ce59",
  1354 => x"e887e6e7",
  1355 => x"d5e787c8",
  1356 => x"c04c7087",
  1357 => x"c102acfb",
  1358 => x"66d487d0",
  1359 => x"87c2c105",
  1360 => x"c11e1ec0",
  1361 => x"faeac11e",
  1362 => x"fd49c01e",
  1363 => x"d0c187eb",
  1364 => x"82c44a66",
  1365 => x"81c7496a",
  1366 => x"1ec15174",
  1367 => x"496a1ed8",
  1368 => x"e5e781c8",
  1369 => x"c186d887",
  1370 => x"c04866c4",
  1371 => x"87c701a8",
  1372 => x"c148a6c4",
  1373 => x"c187ce78",
  1374 => x"c14866c4",
  1375 => x"58a6cc88",
  1376 => x"f1e687c3",
  1377 => x"48a6cc87",
  1378 => x"9c7478c2",
  1379 => x"87cccd02",
  1380 => x"c14866c4",
  1381 => x"03a866c8",
  1382 => x"d887c1cd",
  1383 => x"78c048a6",
  1384 => x"7087e3e5",
  1385 => x"acd0c14c",
  1386 => x"87d6c205",
  1387 => x"e87e66d8",
  1388 => x"497087c7",
  1389 => x"e559a6dc",
  1390 => x"4c7087cc",
  1391 => x"05acecc0",
  1392 => x"c487eac1",
  1393 => x"91cb4966",
  1394 => x"8166c0c1",
  1395 => x"6a4aa1c4",
  1396 => x"4aa1c84d",
  1397 => x"c15266d8",
  1398 => x"e479cfce",
  1399 => x"4c7087e8",
  1400 => x"87d8029c",
  1401 => x"02acfbc0",
  1402 => x"557487d2",
  1403 => x"7087d7e4",
  1404 => x"c7029c4c",
  1405 => x"acfbc087",
  1406 => x"87eeff05",
  1407 => x"c255e0c0",
  1408 => x"97c055c1",
  1409 => x"4966d47d",
  1410 => x"db05a96e",
  1411 => x"4866c487",
  1412 => x"04a866c8",
  1413 => x"66c487ca",
  1414 => x"c880c148",
  1415 => x"87c858a6",
  1416 => x"c14866c8",
  1417 => x"58a6cc88",
  1418 => x"7087dbe3",
  1419 => x"acd0c14c",
  1420 => x"d087c805",
  1421 => x"80c14866",
  1422 => x"c158a6d4",
  1423 => x"fd02acd0",
  1424 => x"a6dc87ea",
  1425 => x"7866d448",
  1426 => x"dc4866d8",
  1427 => x"c905a866",
  1428 => x"e0c087dc",
  1429 => x"f0c048a6",
  1430 => x"cc80c478",
  1431 => x"80c47866",
  1432 => x"747e78c0",
  1433 => x"88fbc048",
  1434 => x"58a6f0c0",
  1435 => x"c8029870",
  1436 => x"cb4887d7",
  1437 => x"a6f0c088",
  1438 => x"02987058",
  1439 => x"4887e9c0",
  1440 => x"f0c088c9",
  1441 => x"987058a6",
  1442 => x"87e1c302",
  1443 => x"c088c448",
  1444 => x"7058a6f0",
  1445 => x"87d60298",
  1446 => x"c088c148",
  1447 => x"7058a6f0",
  1448 => x"c8c30298",
  1449 => x"87dbc787",
  1450 => x"48a6e0c0",
  1451 => x"66cc78c0",
  1452 => x"d080c148",
  1453 => x"cde158a6",
  1454 => x"c04c7087",
  1455 => x"d502acec",
  1456 => x"66e0c087",
  1457 => x"c087c602",
  1458 => x"c95ca6e4",
  1459 => x"c0487487",
  1460 => x"e8c088f0",
  1461 => x"ecc058a6",
  1462 => x"87cc02ac",
  1463 => x"7087e7e0",
  1464 => x"acecc04c",
  1465 => x"87f4ff05",
  1466 => x"1e66e0c0",
  1467 => x"1e4966d4",
  1468 => x"1e66ecc0",
  1469 => x"1efaeac1",
  1470 => x"f64966d4",
  1471 => x"1ec087fb",
  1472 => x"66dc1eca",
  1473 => x"c191cb49",
  1474 => x"d88166d8",
  1475 => x"a1c448a6",
  1476 => x"bf66d878",
  1477 => x"87f2e049",
  1478 => x"b7c086d8",
  1479 => x"c7c106a8",
  1480 => x"de1ec187",
  1481 => x"bf66c81e",
  1482 => x"87dee049",
  1483 => x"497086c8",
  1484 => x"8808c048",
  1485 => x"58a6e4c0",
  1486 => x"06a8b7c0",
  1487 => x"c087e9c0",
  1488 => x"dd4866e0",
  1489 => x"df03a8b7",
  1490 => x"49bf6e87",
  1491 => x"8166e0c0",
  1492 => x"6651e0c0",
  1493 => x"6e81c149",
  1494 => x"c1c281bf",
  1495 => x"66e0c051",
  1496 => x"6e81c249",
  1497 => x"51c081bf",
  1498 => x"dcc47ec1",
  1499 => x"87c9e187",
  1500 => x"58a6e4c0",
  1501 => x"c087c2e1",
  1502 => x"c058a6e8",
  1503 => x"c005a8ec",
  1504 => x"e4c087cb",
  1505 => x"e0c048a6",
  1506 => x"c4c07866",
  1507 => x"f5ddff87",
  1508 => x"4966c487",
  1509 => x"c0c191cb",
  1510 => x"80714866",
  1511 => x"4a6e7e70",
  1512 => x"496e82c8",
  1513 => x"e0c081ca",
  1514 => x"e4c05166",
  1515 => x"81c14966",
  1516 => x"8966e0c0",
  1517 => x"307148c1",
  1518 => x"89c14970",
  1519 => x"c47a9771",
  1520 => x"49bff9c0",
  1521 => x"2966e0c0",
  1522 => x"484a6a97",
  1523 => x"f0c09871",
  1524 => x"496e58a6",
  1525 => x"4d6981c4",
  1526 => x"d84866dc",
  1527 => x"c002a866",
  1528 => x"a6d887c8",
  1529 => x"c078c048",
  1530 => x"a6d887c5",
  1531 => x"d878c148",
  1532 => x"e0c01e66",
  1533 => x"ff49751e",
  1534 => x"c887cfdd",
  1535 => x"c04c7086",
  1536 => x"c106acb7",
  1537 => x"857487d4",
  1538 => x"7449e0c0",
  1539 => x"c14b7589",
  1540 => x"714ad4e4",
  1541 => x"87cee3fe",
  1542 => x"e8c085c2",
  1543 => x"80c14866",
  1544 => x"58a6ecc0",
  1545 => x"4966ecc0",
  1546 => x"a97081c1",
  1547 => x"87c8c002",
  1548 => x"c048a6d8",
  1549 => x"87c5c078",
  1550 => x"c148a6d8",
  1551 => x"1e66d878",
  1552 => x"c049a4c2",
  1553 => x"887148e0",
  1554 => x"751e4970",
  1555 => x"f9dbff49",
  1556 => x"c086c887",
  1557 => x"ff01a8b7",
  1558 => x"e8c087c0",
  1559 => x"d1c00266",
  1560 => x"c9496e87",
  1561 => x"66e8c081",
  1562 => x"c1486e51",
  1563 => x"c078dfcf",
  1564 => x"496e87cc",
  1565 => x"51c281c9",
  1566 => x"d0c1486e",
  1567 => x"7ec178d3",
  1568 => x"ff87c6c0",
  1569 => x"7087efda",
  1570 => x"c0026e4c",
  1571 => x"66c487f5",
  1572 => x"a866c848",
  1573 => x"87cbc004",
  1574 => x"c14866c4",
  1575 => x"58a6c880",
  1576 => x"c887e0c0",
  1577 => x"88c14866",
  1578 => x"c058a6cc",
  1579 => x"c6c187d5",
  1580 => x"c8c005ac",
  1581 => x"4866cc87",
  1582 => x"a6d080c1",
  1583 => x"f5d9ff58",
  1584 => x"d04c7087",
  1585 => x"80c14866",
  1586 => x"7458a6d4",
  1587 => x"cbc0029c",
  1588 => x"4866c487",
  1589 => x"a866c8c1",
  1590 => x"87fff204",
  1591 => x"87cdd9ff",
  1592 => x"c74866c4",
  1593 => x"e5c003a8",
  1594 => x"ccfdc387",
  1595 => x"c478c048",
  1596 => x"91cb4966",
  1597 => x"8166c0c1",
  1598 => x"6a4aa1c4",
  1599 => x"7952c04a",
  1600 => x"c14866c4",
  1601 => x"58a6c880",
  1602 => x"ff04a8c7",
  1603 => x"d0ff87db",
  1604 => x"87f5e08e",
  1605 => x"1e00203a",
  1606 => x"4b711e73",
  1607 => x"87c6029b",
  1608 => x"48c8fdc3",
  1609 => x"1ec778c0",
  1610 => x"bfc8fdc3",
  1611 => x"e9c11e49",
  1612 => x"fdc31ed7",
  1613 => x"ee49bfc4",
  1614 => x"86cc87f4",
  1615 => x"bfc4fdc3",
  1616 => x"87f3e949",
  1617 => x"c8029b73",
  1618 => x"d7e9c187",
  1619 => x"c2e7c049",
  1620 => x"f8dfff87",
  1621 => x"1e731e87",
  1622 => x"4bffc31e",
  1623 => x"fc4ad4ff",
  1624 => x"98c148bf",
  1625 => x"026e7e70",
  1626 => x"ff87fbc0",
  1627 => x"c1c148d0",
  1628 => x"7ad2c278",
  1629 => x"f0c37a73",
  1630 => x"ff4849d3",
  1631 => x"73506a80",
  1632 => x"73516a7a",
  1633 => x"6a80c17a",
  1634 => x"6a7a7350",
  1635 => x"6a7a7350",
  1636 => x"6a7a7349",
  1637 => x"6a7a7350",
  1638 => x"dcf0c350",
  1639 => x"d0ff5997",
  1640 => x"78c0c148",
  1641 => x"f0c387d7",
  1642 => x"ff4849d3",
  1643 => x"5150c080",
  1644 => x"50c080c1",
  1645 => x"50c150d9",
  1646 => x"c350e2c0",
  1647 => x"d9f0c350",
  1648 => x"f850c048",
  1649 => x"deff2680",
  1650 => x"c71e87c3",
  1651 => x"49c187cb",
  1652 => x"fe87c4fd",
  1653 => x"7087d4e6",
  1654 => x"87cd0298",
  1655 => x"87d1effe",
  1656 => x"c4029870",
  1657 => x"c24ac187",
  1658 => x"724ac087",
  1659 => x"87ce059a",
  1660 => x"e8c11ec0",
  1661 => x"f0c049db",
  1662 => x"86c487f4",
  1663 => x"1ec087fe",
  1664 => x"49e6e8c1",
  1665 => x"87e6f0c0",
  1666 => x"fbc11ec0",
  1667 => x"497087c6",
  1668 => x"87daf0c0",
  1669 => x"f887c1c3",
  1670 => x"534f268e",
  1671 => x"61662044",
  1672 => x"64656c69",
  1673 => x"6f42002e",
  1674 => x"6e69746f",
  1675 => x"2e2e2e67",
  1676 => x"fdc31e00",
  1677 => x"78c048c8",
  1678 => x"48c4fdc3",
  1679 => x"c9fe78c0",
  1680 => x"f6fdc187",
  1681 => x"2648c087",
  1682 => x"4520804f",
  1683 => x"00746978",
  1684 => x"61422080",
  1685 => x"8f006b63",
  1686 => x"5d000013",
  1687 => x"0000003f",
  1688 => x"138f0000",
  1689 => x"3f7b0000",
  1690 => x"00000000",
  1691 => x"00138f00",
  1692 => x"003f9900",
  1693 => x"00000000",
  1694 => x"0000138f",
  1695 => x"00003fb7",
  1696 => x"8f000000",
  1697 => x"d5000013",
  1698 => x"0000003f",
  1699 => x"138f0000",
  1700 => x"3ff30000",
  1701 => x"00000000",
  1702 => x"00138f00",
  1703 => x"00401100",
  1704 => x"00000000",
  1705 => x"0000138f",
  1706 => x"00000000",
  1707 => x"2a000000",
  1708 => x"00000014",
  1709 => x"00000000",
  1710 => x"6f4c0000",
  1711 => x"2a206461",
  1712 => x"fe1e002e",
  1713 => x"78c048f0",
  1714 => x"097909cd",
  1715 => x"1e1e4f26",
  1716 => x"7ebff0fe",
  1717 => x"4f262648",
  1718 => x"48f0fe1e",
  1719 => x"4f2678c1",
  1720 => x"48f0fe1e",
  1721 => x"4f2678c0",
  1722 => x"c04a711e",
  1723 => x"4f265252",
  1724 => x"5c5b5e0e",
  1725 => x"86f40e5d",
  1726 => x"6d974d71",
  1727 => x"4ca5c17e",
  1728 => x"c8486c97",
  1729 => x"486e58a6",
  1730 => x"05a866c4",
  1731 => x"48ff87c5",
  1732 => x"ff87e6c0",
  1733 => x"a5c287ca",
  1734 => x"4b6c9749",
  1735 => x"974ba371",
  1736 => x"6c974b6b",
  1737 => x"c1486e7e",
  1738 => x"58a6c880",
  1739 => x"a6cc98c7",
  1740 => x"7c977058",
  1741 => x"7387e1fe",
  1742 => x"268ef448",
  1743 => x"264c264d",
  1744 => x"0e4f264b",
  1745 => x"0e5c5b5e",
  1746 => x"4c7186f4",
  1747 => x"c34a66d8",
  1748 => x"a4c29aff",
  1749 => x"496c974b",
  1750 => x"7249a173",
  1751 => x"7e6c9751",
  1752 => x"80c1486e",
  1753 => x"c758a6c8",
  1754 => x"58a6cc98",
  1755 => x"8ef45470",
  1756 => x"1e87caff",
  1757 => x"87e8fd1e",
  1758 => x"494abfe0",
  1759 => x"99c0e0c0",
  1760 => x"7287cb02",
  1761 => x"efc0c41e",
  1762 => x"87f7fe49",
  1763 => x"fdfc86c4",
  1764 => x"fd7e7087",
  1765 => x"262687c2",
  1766 => x"c0c41e4f",
  1767 => x"c7fd49ef",
  1768 => x"f3edc187",
  1769 => x"87dafc49",
  1770 => x"2687f8c4",
  1771 => x"5b5e0e4f",
  1772 => x"c40e5d5c",
  1773 => x"4abfcec1",
  1774 => x"bfc1f0c1",
  1775 => x"bc724c49",
  1776 => x"dbfc4d71",
  1777 => x"744bc087",
  1778 => x"0299d049",
  1779 => x"497587d5",
  1780 => x"1e7199d0",
  1781 => x"f5c11ec0",
  1782 => x"82734af2",
  1783 => x"e4c04912",
  1784 => x"c186c887",
  1785 => x"c8832d2c",
  1786 => x"daff04ab",
  1787 => x"87e8fb87",
  1788 => x"48c1f0c1",
  1789 => x"bfcec1c4",
  1790 => x"264d2678",
  1791 => x"264b264c",
  1792 => x"0000004f",
  1793 => x"d0ff1e00",
  1794 => x"78e1c848",
  1795 => x"c548d4ff",
  1796 => x"0266c478",
  1797 => x"e0c387c3",
  1798 => x"0266c878",
  1799 => x"d4ff87c6",
  1800 => x"78f0c348",
  1801 => x"7148d4ff",
  1802 => x"48d0ff78",
  1803 => x"c078e1c8",
  1804 => x"4f2678e0",
  1805 => x"c41e731e",
  1806 => x"fa49efc0",
  1807 => x"4a7087f2",
  1808 => x"04aab7c0",
  1809 => x"c387cfc2",
  1810 => x"c905aae0",
  1811 => x"dff3c187",
  1812 => x"c278c148",
  1813 => x"497287c0",
  1814 => x"0299c0c2",
  1815 => x"f3c187c9",
  1816 => x"78c148db",
  1817 => x"c19afffd",
  1818 => x"02bfdff3",
  1819 => x"4b7287c7",
  1820 => x"c2b3c0c2",
  1821 => x"c14b7287",
  1822 => x"02bfdbf3",
  1823 => x"7387e0c0",
  1824 => x"29b7c449",
  1825 => x"f2f4c191",
  1826 => x"cf4a7381",
  1827 => x"c192c29a",
  1828 => x"70307248",
  1829 => x"72baff4a",
  1830 => x"70986948",
  1831 => x"7387db79",
  1832 => x"29b7c449",
  1833 => x"f2f4c191",
  1834 => x"cf4a7381",
  1835 => x"c392c29a",
  1836 => x"70307248",
  1837 => x"b069484a",
  1838 => x"f3c17970",
  1839 => x"78c048df",
  1840 => x"48dbf3c1",
  1841 => x"c0c478c0",
  1842 => x"e3f849ef",
  1843 => x"c04a7087",
  1844 => x"fd03aab7",
  1845 => x"48c087f1",
  1846 => x"0087e2fc",
  1847 => x"00000000",
  1848 => x"1e000000",
  1849 => x"49724ac0",
  1850 => x"f4c191c4",
  1851 => x"79c081f2",
  1852 => x"b7d082c1",
  1853 => x"87ee04aa",
  1854 => x"5e0e4f26",
  1855 => x"0e5d5c5b",
  1856 => x"dbf74d71",
  1857 => x"c44a7587",
  1858 => x"c1922ab7",
  1859 => x"7582f2f4",
  1860 => x"c29ccf4c",
  1861 => x"4b496a94",
  1862 => x"9bc32b74",
  1863 => x"307448c2",
  1864 => x"bcff4c70",
  1865 => x"98714874",
  1866 => x"ebf67a70",
  1867 => x"fb487387",
  1868 => x"000087c7",
  1869 => x"00000000",
  1870 => x"00000000",
  1871 => x"00000000",
  1872 => x"00000000",
  1873 => x"00000000",
  1874 => x"00000000",
  1875 => x"00000000",
  1876 => x"00000000",
  1877 => x"00000000",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"00000000",
  1884 => x"1e160000",
  1885 => x"362e2526",
  1886 => x"ff1e3e3d",
  1887 => x"e1c848d0",
  1888 => x"ff487178",
  1889 => x"267808d4",
  1890 => x"d0ff1e4f",
  1891 => x"78e1c848",
  1892 => x"d4ff4871",
  1893 => x"66c47808",
  1894 => x"08d4ff48",
  1895 => x"1e4f2678",
  1896 => x"66c44a71",
  1897 => x"49721e49",
  1898 => x"ff87deff",
  1899 => x"e0c048d0",
  1900 => x"4f262678",
  1901 => x"c44a711e",
  1902 => x"e0c11e66",
  1903 => x"c8ff49a2",
  1904 => x"4966c887",
  1905 => x"ff29b7c8",
  1906 => x"787148d4",
  1907 => x"c048d0ff",
  1908 => x"262678e0",
  1909 => x"1e731e4f",
  1910 => x"e2c04b71",
  1911 => x"87dafe49",
  1912 => x"48134ac7",
  1913 => x"7808d4ff",
  1914 => x"8ac14972",
  1915 => x"f1059971",
  1916 => x"48d0ff87",
  1917 => x"c478e0c0",
  1918 => x"264d2687",
  1919 => x"264b264c",
  1920 => x"d4ff1e4f",
  1921 => x"7affc34a",
  1922 => x"c848d0ff",
  1923 => x"7ade78e1",
  1924 => x"bff9c0c4",
  1925 => x"c848497a",
  1926 => x"717a7028",
  1927 => x"7028d048",
  1928 => x"d848717a",
  1929 => x"ff7a7028",
  1930 => x"e0c048d0",
  1931 => x"0e4f2678",
  1932 => x"5d5c5b5e",
  1933 => x"c44c710e",
  1934 => x"4dbff9c0",
  1935 => x"d02b744b",
  1936 => x"83c19b66",
  1937 => x"04ab66d4",
  1938 => x"4bc087c2",
  1939 => x"66d04a74",
  1940 => x"ff317249",
  1941 => x"739975b9",
  1942 => x"70307248",
  1943 => x"b071484a",
  1944 => x"58fdc0c4",
  1945 => x"2687dafe",
  1946 => x"264c264d",
  1947 => x"1e4f264b",
  1948 => x"c848d0ff",
  1949 => x"487178c9",
  1950 => x"7808d4ff",
  1951 => x"711e4f26",
  1952 => x"87eb494a",
  1953 => x"c848d0ff",
  1954 => x"1e4f2678",
  1955 => x"4b711e73",
  1956 => x"bfc9c1c4",
  1957 => x"c287c302",
  1958 => x"d0ff87eb",
  1959 => x"78c9c848",
  1960 => x"e0c04973",
  1961 => x"48d4ffb1",
  1962 => x"c0c47871",
  1963 => x"78c048fd",
  1964 => x"c50266c8",
  1965 => x"49ffc387",
  1966 => x"49c087c2",
  1967 => x"59c5c1c4",
  1968 => x"c60266cc",
  1969 => x"d5d5c587",
  1970 => x"cf87c44a",
  1971 => x"c44affff",
  1972 => x"c45ac9c1",
  1973 => x"c148c9c1",
  1974 => x"2687c478",
  1975 => x"264c264d",
  1976 => x"0e4f264b",
  1977 => x"5d5c5b5e",
  1978 => x"c44a710e",
  1979 => x"4cbfc5c1",
  1980 => x"cb029a72",
  1981 => x"91c84987",
  1982 => x"4bc1fac1",
  1983 => x"87c48371",
  1984 => x"4bc1fec1",
  1985 => x"49134dc0",
  1986 => x"c1c49974",
  1987 => x"ffb9bfc1",
  1988 => x"787148d4",
  1989 => x"852cb7c1",
  1990 => x"04adb7c8",
  1991 => x"c0c487e8",
  1992 => x"c848bffd",
  1993 => x"c1c1c480",
  1994 => x"87effe58",
  1995 => x"711e731e",
  1996 => x"9a4a134b",
  1997 => x"7287cb02",
  1998 => x"87e7fe49",
  1999 => x"059a4a13",
  2000 => x"dafe87f5",
  2001 => x"c0c41e87",
  2002 => x"c449bffd",
  2003 => x"c148fdc0",
  2004 => x"c0c478a1",
  2005 => x"db03a9b7",
  2006 => x"48d4ff87",
  2007 => x"bfc1c1c4",
  2008 => x"fdc0c478",
  2009 => x"c0c449bf",
  2010 => x"a1c148fd",
  2011 => x"b7c0c478",
  2012 => x"87e504a9",
  2013 => x"c848d0ff",
  2014 => x"c9c1c478",
  2015 => x"2678c048",
  2016 => x"0000004f",
  2017 => x"00000000",
  2018 => x"00000000",
  2019 => x"00005f5f",
  2020 => x"03030000",
  2021 => x"00030300",
  2022 => x"7f7f1400",
  2023 => x"147f7f14",
  2024 => x"2e240000",
  2025 => x"123a6b6b",
  2026 => x"366a4c00",
  2027 => x"32566c18",
  2028 => x"4f7e3000",
  2029 => x"683a7759",
  2030 => x"04000040",
  2031 => x"00000307",
  2032 => x"1c000000",
  2033 => x"0041633e",
  2034 => x"41000000",
  2035 => x"001c3e63",
  2036 => x"3e2a0800",
  2037 => x"2a3e1c1c",
  2038 => x"08080008",
  2039 => x"08083e3e",
  2040 => x"80000000",
  2041 => x"000060e0",
  2042 => x"08080000",
  2043 => x"08080808",
  2044 => x"00000000",
  2045 => x"00006060",
  2046 => x"30604000",
  2047 => x"03060c18",
  2048 => x"7f3e0001",
  2049 => x"3e7f4d59",
  2050 => x"06040000",
  2051 => x"00007f7f",
  2052 => x"63420000",
  2053 => x"464f5971",
  2054 => x"63220000",
  2055 => x"367f4949",
  2056 => x"161c1800",
  2057 => x"107f7f13",
  2058 => x"67270000",
  2059 => x"397d4545",
  2060 => x"7e3c0000",
  2061 => x"3079494b",
  2062 => x"01010000",
  2063 => x"070f7971",
  2064 => x"7f360000",
  2065 => x"367f4949",
  2066 => x"4f060000",
  2067 => x"1e3f6949",
  2068 => x"00000000",
  2069 => x"00006666",
  2070 => x"80000000",
  2071 => x"000066e6",
  2072 => x"08080000",
  2073 => x"22221414",
  2074 => x"14140000",
  2075 => x"14141414",
  2076 => x"22220000",
  2077 => x"08081414",
  2078 => x"03020000",
  2079 => x"060f5951",
  2080 => x"417f3e00",
  2081 => x"1e1f555d",
  2082 => x"7f7e0000",
  2083 => x"7e7f0909",
  2084 => x"7f7f0000",
  2085 => x"367f4949",
  2086 => x"3e1c0000",
  2087 => x"41414163",
  2088 => x"7f7f0000",
  2089 => x"1c3e6341",
  2090 => x"7f7f0000",
  2091 => x"41414949",
  2092 => x"7f7f0000",
  2093 => x"01010909",
  2094 => x"7f3e0000",
  2095 => x"7a7b4941",
  2096 => x"7f7f0000",
  2097 => x"7f7f0808",
  2098 => x"41000000",
  2099 => x"00417f7f",
  2100 => x"60200000",
  2101 => x"3f7f4040",
  2102 => x"087f7f00",
  2103 => x"4163361c",
  2104 => x"7f7f0000",
  2105 => x"40404040",
  2106 => x"067f7f00",
  2107 => x"7f7f060c",
  2108 => x"067f7f00",
  2109 => x"7f7f180c",
  2110 => x"7f3e0000",
  2111 => x"3e7f4141",
  2112 => x"7f7f0000",
  2113 => x"060f0909",
  2114 => x"417f3e00",
  2115 => x"407e7f61",
  2116 => x"7f7f0000",
  2117 => x"667f1909",
  2118 => x"6f260000",
  2119 => x"327b594d",
  2120 => x"01010000",
  2121 => x"01017f7f",
  2122 => x"7f3f0000",
  2123 => x"3f7f4040",
  2124 => x"3f0f0000",
  2125 => x"0f3f7070",
  2126 => x"307f7f00",
  2127 => x"7f7f3018",
  2128 => x"36634100",
  2129 => x"63361c1c",
  2130 => x"06030141",
  2131 => x"03067c7c",
  2132 => x"59716101",
  2133 => x"4143474d",
  2134 => x"7f000000",
  2135 => x"0041417f",
  2136 => x"06030100",
  2137 => x"6030180c",
  2138 => x"41000040",
  2139 => x"007f7f41",
  2140 => x"060c0800",
  2141 => x"080c0603",
  2142 => x"80808000",
  2143 => x"80808080",
  2144 => x"00000000",
  2145 => x"00040703",
  2146 => x"74200000",
  2147 => x"787c5454",
  2148 => x"7f7f0000",
  2149 => x"387c4444",
  2150 => x"7c380000",
  2151 => x"00444444",
  2152 => x"7c380000",
  2153 => x"7f7f4444",
  2154 => x"7c380000",
  2155 => x"185c5454",
  2156 => x"7e040000",
  2157 => x"0005057f",
  2158 => x"bc180000",
  2159 => x"7cfca4a4",
  2160 => x"7f7f0000",
  2161 => x"787c0404",
  2162 => x"00000000",
  2163 => x"00407d3d",
  2164 => x"80800000",
  2165 => x"007dfd80",
  2166 => x"7f7f0000",
  2167 => x"446c3810",
  2168 => x"00000000",
  2169 => x"00407f3f",
  2170 => x"0c7c7c00",
  2171 => x"787c0c18",
  2172 => x"7c7c0000",
  2173 => x"787c0404",
  2174 => x"7c380000",
  2175 => x"387c4444",
  2176 => x"fcfc0000",
  2177 => x"183c2424",
  2178 => x"3c180000",
  2179 => x"fcfc2424",
  2180 => x"7c7c0000",
  2181 => x"080c0404",
  2182 => x"5c480000",
  2183 => x"20745454",
  2184 => x"3f040000",
  2185 => x"0044447f",
  2186 => x"7c3c0000",
  2187 => x"7c7c4040",
  2188 => x"3c1c0000",
  2189 => x"1c3c6060",
  2190 => x"607c3c00",
  2191 => x"3c7c6030",
  2192 => x"386c4400",
  2193 => x"446c3810",
  2194 => x"bc1c0000",
  2195 => x"1c3c60e0",
  2196 => x"64440000",
  2197 => x"444c5c74",
  2198 => x"08080000",
  2199 => x"4141773e",
  2200 => x"00000000",
  2201 => x"00007f7f",
  2202 => x"41410000",
  2203 => x"08083e77",
  2204 => x"01010200",
  2205 => x"01020203",
  2206 => x"7f7f7f00",
  2207 => x"7f7f7f7f",
  2208 => x"1c080800",
  2209 => x"7f3e3e1c",
  2210 => x"3e7f7f7f",
  2211 => x"081c1c3e",
  2212 => x"18100008",
  2213 => x"10187c7c",
  2214 => x"30100000",
  2215 => x"10307c7c",
  2216 => x"60301000",
  2217 => x"061e7860",
  2218 => x"3c664200",
  2219 => x"42663c18",
  2220 => x"6a387800",
  2221 => x"386cc6c2",
  2222 => x"00006000",
  2223 => x"60000060",
  2224 => x"5b5e0e00",
  2225 => x"1e0e5d5c",
  2226 => x"c1c44c71",
  2227 => x"c04dbfda",
  2228 => x"741ec04b",
  2229 => x"87c702ab",
  2230 => x"c048a6c4",
  2231 => x"c487c578",
  2232 => x"78c148a6",
  2233 => x"731e66c4",
  2234 => x"87dfee49",
  2235 => x"e0c086c8",
  2236 => x"87efef49",
  2237 => x"6a4aa5c4",
  2238 => x"87f0f049",
  2239 => x"cb87c6f1",
  2240 => x"c883c185",
  2241 => x"ff04abb7",
  2242 => x"262687c7",
  2243 => x"264c264d",
  2244 => x"1e4f264b",
  2245 => x"c1c44a71",
  2246 => x"c1c45ade",
  2247 => x"78c748de",
  2248 => x"87ddfe49",
  2249 => x"731e4f26",
  2250 => x"c04a711e",
  2251 => x"d303aab7",
  2252 => x"c3dac287",
  2253 => x"87c405bf",
  2254 => x"87c24bc1",
  2255 => x"dac24bc0",
  2256 => x"87c45bc7",
  2257 => x"5ac7dac2",
  2258 => x"bfc3dac2",
  2259 => x"c19ac14a",
  2260 => x"ec49a2c0",
  2261 => x"48fc87e8",
  2262 => x"bfc3dac2",
  2263 => x"87effe78",
  2264 => x"c3dac21e",
  2265 => x"4f2648bf",
  2266 => x"c44a711e",
  2267 => x"49721e66",
  2268 => x"2687c1e9",
  2269 => x"c21e4f26",
  2270 => x"49bfc3da",
  2271 => x"87dcd2c1",
  2272 => x"48d2c1c4",
  2273 => x"c478bfe8",
  2274 => x"ec48cec1",
  2275 => x"c1c478bf",
  2276 => x"494abfd2",
  2277 => x"c899ffc3",
  2278 => x"48722ab7",
  2279 => x"c1c4b071",
  2280 => x"4f2658da",
  2281 => x"5c5b5e0e",
  2282 => x"4b710e5d",
  2283 => x"c487c7ff",
  2284 => x"c048cdc1",
  2285 => x"e5497350",
  2286 => x"497087c0",
  2287 => x"cb9cc24c",
  2288 => x"c6cb49ee",
  2289 => x"4d497087",
  2290 => x"97cdc1c4",
  2291 => x"e2c105bf",
  2292 => x"4966d087",
  2293 => x"bfd6c1c4",
  2294 => x"87d60599",
  2295 => x"c44966d4",
  2296 => x"99bfcec1",
  2297 => x"7387cb05",
  2298 => x"87cee449",
  2299 => x"c1029870",
  2300 => x"4cc187c1",
  2301 => x"7587fffd",
  2302 => x"87dbca49",
  2303 => x"c6029870",
  2304 => x"cdc1c487",
  2305 => x"c450c148",
  2306 => x"bf97cdc1",
  2307 => x"87e3c005",
  2308 => x"bfd6c1c4",
  2309 => x"9966d049",
  2310 => x"87d6ff05",
  2311 => x"bfcec1c4",
  2312 => x"9966d449",
  2313 => x"87caff05",
  2314 => x"cde34973",
  2315 => x"05987087",
  2316 => x"7487fffe",
  2317 => x"87d3fb48",
  2318 => x"5c5b5e0e",
  2319 => x"86f40e5d",
  2320 => x"ec4c4dc0",
  2321 => x"a6c47ebf",
  2322 => x"dac1c448",
  2323 => x"1ec178bf",
  2324 => x"d8c11ec0",
  2325 => x"87ccfd49",
  2326 => x"987086c8",
  2327 => x"ff87cc02",
  2328 => x"87c2fb49",
  2329 => x"d1e249dc",
  2330 => x"c44dc187",
  2331 => x"bf97cdc1",
  2332 => x"c087c402",
  2333 => x"c487e4fd",
  2334 => x"4bbfd2c1",
  2335 => x"bfc3dac2",
  2336 => x"87e9c005",
  2337 => x"e149c9c3",
  2338 => x"e1c387f0",
  2339 => x"87eae149",
  2340 => x"ffc34973",
  2341 => x"c01e7199",
  2342 => x"87ccfb49",
  2343 => x"b7c84973",
  2344 => x"c11e7129",
  2345 => x"87c0fb49",
  2346 => x"fcc586c8",
  2347 => x"d6c1c487",
  2348 => x"029b4bbf",
  2349 => x"d9c287dd",
  2350 => x"c749bfff",
  2351 => x"987087d9",
  2352 => x"c087c405",
  2353 => x"c287d24b",
  2354 => x"fec649e0",
  2355 => x"c3dac287",
  2356 => x"c287c658",
  2357 => x"c048ffd9",
  2358 => x"c2497378",
  2359 => x"87cd0599",
  2360 => x"e049cbc3",
  2361 => x"497087d4",
  2362 => x"c20299c2",
  2363 => x"734cfb87",
  2364 => x"0599c149",
  2365 => x"cdc387ce",
  2366 => x"fddfff49",
  2367 => x"c2497087",
  2368 => x"87c20299",
  2369 => x"49734cfa",
  2370 => x"ce0599c8",
  2371 => x"49c8c387",
  2372 => x"87e6dfff",
  2373 => x"99c24970",
  2374 => x"c487d502",
  2375 => x"02bfdec1",
  2376 => x"c14887ca",
  2377 => x"e2c1c488",
  2378 => x"87c2c058",
  2379 => x"4dc14cff",
  2380 => x"99c44973",
  2381 => x"c387ce05",
  2382 => x"deff49d0",
  2383 => x"497087fc",
  2384 => x"db0299c2",
  2385 => x"dec1c487",
  2386 => x"c7487ebf",
  2387 => x"cb03a8b7",
  2388 => x"c1486e87",
  2389 => x"e2c1c480",
  2390 => x"87c2c058",
  2391 => x"4dc14cfe",
  2392 => x"ff49c9c3",
  2393 => x"7087d3de",
  2394 => x"0299c249",
  2395 => x"c1c487d5",
  2396 => x"c002bfde",
  2397 => x"c1c487c9",
  2398 => x"78c048de",
  2399 => x"fd87c2c0",
  2400 => x"c34dc14c",
  2401 => x"ddff49e1",
  2402 => x"497087f0",
  2403 => x"d90299c2",
  2404 => x"dec1c487",
  2405 => x"b7c748bf",
  2406 => x"c9c003a8",
  2407 => x"dec1c487",
  2408 => x"c078c748",
  2409 => x"4cfc87c2",
  2410 => x"b7c04dc1",
  2411 => x"d1c003ac",
  2412 => x"4a66c487",
  2413 => x"6a82d8c1",
  2414 => x"87c6c002",
  2415 => x"49744b6a",
  2416 => x"1ec00f73",
  2417 => x"dc1ef0c3",
  2418 => x"87d8f749",
  2419 => x"987086c8",
  2420 => x"87e2c002",
  2421 => x"c448a6c8",
  2422 => x"78bfdec1",
  2423 => x"cb4966c8",
  2424 => x"4866c491",
  2425 => x"7e708071",
  2426 => x"c002bf6e",
  2427 => x"bf6e87c8",
  2428 => x"4966c84b",
  2429 => x"9d750f73",
  2430 => x"87c8c002",
  2431 => x"bfdec1c4",
  2432 => x"87fdf249",
  2433 => x"bfc7dac2",
  2434 => x"87ddc002",
  2435 => x"87c7c249",
  2436 => x"c0029870",
  2437 => x"c1c487d3",
  2438 => x"f249bfde",
  2439 => x"49c087e3",
  2440 => x"c287c3f4",
  2441 => x"c048c7da",
  2442 => x"f38ef478",
  2443 => x"5e0e87dd",
  2444 => x"0e5d5c5b",
  2445 => x"c44c711e",
  2446 => x"49bfdac1",
  2447 => x"4da1cdc1",
  2448 => x"6981d1c1",
  2449 => x"029c747e",
  2450 => x"a5c487cf",
  2451 => x"c47b744b",
  2452 => x"49bfdac1",
  2453 => x"6e87fcf2",
  2454 => x"059c747b",
  2455 => x"4bc087c4",
  2456 => x"4bc187c2",
  2457 => x"fdf24973",
  2458 => x"0266d487",
  2459 => x"da4987c7",
  2460 => x"c24a7087",
  2461 => x"c24ac087",
  2462 => x"265acbda",
  2463 => x"0087ccf2",
  2464 => x"00000000",
  2465 => x"00000000",
  2466 => x"1e000000",
  2467 => x"c8ff4a71",
  2468 => x"a17249bf",
  2469 => x"1e4f2648",
  2470 => x"89bfc8ff",
  2471 => x"c0c0c0fe",
  2472 => x"01a9c0c0",
  2473 => x"4ac087c4",
  2474 => x"4ac187c2",
  2475 => x"4f264872",
  2476 => x"5c5b5e0e",
  2477 => x"4b710e5d",
  2478 => x"d04cd4ff",
  2479 => x"78c04866",
  2480 => x"daff49d6",
  2481 => x"ffc387f4",
  2482 => x"c3496c7c",
  2483 => x"4d7199ff",
  2484 => x"99f0c349",
  2485 => x"05a9e0c1",
  2486 => x"ffc387cb",
  2487 => x"c3486c7c",
  2488 => x"0866d098",
  2489 => x"7cffc378",
  2490 => x"c8494a6c",
  2491 => x"7cffc331",
  2492 => x"b2714a6c",
  2493 => x"31c84972",
  2494 => x"6c7cffc3",
  2495 => x"72b2714a",
  2496 => x"c331c849",
  2497 => x"4a6c7cff",
  2498 => x"d0ffb271",
  2499 => x"78e0c048",
  2500 => x"c2029b73",
  2501 => x"757b7287",
  2502 => x"264d2648",
  2503 => x"264b264c",
  2504 => x"4f261e4f",
  2505 => x"5c5b5e0e",
  2506 => x"7686f80e",
  2507 => x"49a6c81e",
  2508 => x"c487fdfd",
  2509 => x"6e4b7086",
  2510 => x"03a8c248",
  2511 => x"7387cac3",
  2512 => x"9af0c34a",
  2513 => x"02aad0c1",
  2514 => x"e0c187c7",
  2515 => x"f8c205aa",
  2516 => x"c8497387",
  2517 => x"87c30299",
  2518 => x"7387c6ff",
  2519 => x"c29cc34c",
  2520 => x"cfc105ac",
  2521 => x"4966c487",
  2522 => x"1e7131c9",
  2523 => x"c24a66c4",
  2524 => x"c1c492d8",
  2525 => x"817249e2",
  2526 => x"87c2d0fe",
  2527 => x"1e4966c4",
  2528 => x"ff49e3c0",
  2529 => x"d887d8d8",
  2530 => x"edd7ff49",
  2531 => x"1ec0c887",
  2532 => x"49d2f0c3",
  2533 => x"87f3e7fd",
  2534 => x"c048d0ff",
  2535 => x"f0c378e0",
  2536 => x"66d01ed2",
  2537 => x"92d8c24a",
  2538 => x"49e2c1c4",
  2539 => x"cafe8172",
  2540 => x"86d087dd",
  2541 => x"c105acc1",
  2542 => x"66c487cf",
  2543 => x"7131c949",
  2544 => x"4a66c41e",
  2545 => x"c492d8c2",
  2546 => x"7249e2c1",
  2547 => x"edcefe81",
  2548 => x"d2f0c387",
  2549 => x"4a66c81e",
  2550 => x"c492d8c2",
  2551 => x"7249e2c1",
  2552 => x"e7c8fe81",
  2553 => x"4966c887",
  2554 => x"49e3c01e",
  2555 => x"87efd6ff",
  2556 => x"d6ff49d7",
  2557 => x"c0c887c4",
  2558 => x"d2f0c31e",
  2559 => x"f4e5fd49",
  2560 => x"ff86d087",
  2561 => x"e0c048d0",
  2562 => x"fc8ef878",
  2563 => x"5e0e87cd",
  2564 => x"0e5d5c5b",
  2565 => x"ff4d711e",
  2566 => x"66d44cd4",
  2567 => x"b7c3487e",
  2568 => x"87c506a8",
  2569 => x"e3c148c0",
  2570 => x"fe497587",
  2571 => x"7587f7df",
  2572 => x"4b66c41e",
  2573 => x"c493d8c2",
  2574 => x"7383e2c1",
  2575 => x"fec2fe49",
  2576 => x"6b83c887",
  2577 => x"48d0ff4b",
  2578 => x"dd78e1c8",
  2579 => x"c349737c",
  2580 => x"7c7199ff",
  2581 => x"b7c84973",
  2582 => x"99ffc329",
  2583 => x"49737c71",
  2584 => x"c329b7d0",
  2585 => x"7c7199ff",
  2586 => x"b7d84973",
  2587 => x"c07c7129",
  2588 => x"7c7c7c7c",
  2589 => x"7c7c7c7c",
  2590 => x"7c7c7c7c",
  2591 => x"c478e0c0",
  2592 => x"49dc1e66",
  2593 => x"87d7d4ff",
  2594 => x"487386c8",
  2595 => x"87c9fa26",
  2596 => x"4ad4ff1e",
  2597 => x"c848d0ff",
  2598 => x"f0c378c5",
  2599 => x"c07a717a",
  2600 => x"7a7a7a7a",
  2601 => x"4f2678c4",
  2602 => x"4ad4ff1e",
  2603 => x"c848d0ff",
  2604 => x"7ac078c5",
  2605 => x"7ac0496a",
  2606 => x"7a7a7a7a",
  2607 => x"487178c4",
  2608 => x"5e0e4f26",
  2609 => x"0e5d5c5b",
  2610 => x"a6cc86e4",
  2611 => x"66ecc059",
  2612 => x"58a6dc48",
  2613 => x"e8c24d70",
  2614 => x"d2c6c495",
  2615 => x"a5d8c285",
  2616 => x"48a6c47e",
  2617 => x"78a5dcc2",
  2618 => x"4cbf66c4",
  2619 => x"c294bf6e",
  2620 => x"946d85e0",
  2621 => x"c04b66c8",
  2622 => x"49c0c84a",
  2623 => x"87c3e0fd",
  2624 => x"c14866c8",
  2625 => x"c8789fc0",
  2626 => x"81c24966",
  2627 => x"799fbf6e",
  2628 => x"c64966c8",
  2629 => x"bf66c481",
  2630 => x"66c8799f",
  2631 => x"6d81cc49",
  2632 => x"66c8799f",
  2633 => x"d080d448",
  2634 => x"e7c258a6",
  2635 => x"66cc48fb",
  2636 => x"4aa1d449",
  2637 => x"aa714120",
  2638 => x"c887f905",
  2639 => x"eec04866",
  2640 => x"58a6d480",
  2641 => x"48d0e8c2",
  2642 => x"c84966d0",
  2643 => x"41204aa1",
  2644 => x"f905aa71",
  2645 => x"4866c887",
  2646 => x"d880f6c0",
  2647 => x"e8c258a6",
  2648 => x"66d448d9",
  2649 => x"a1e8c049",
  2650 => x"7141204a",
  2651 => x"87f905aa",
  2652 => x"c04a66d8",
  2653 => x"66d482f1",
  2654 => x"7281cb49",
  2655 => x"4966c851",
  2656 => x"c881dec1",
  2657 => x"799fd0c0",
  2658 => x"c14966c8",
  2659 => x"c0c881e2",
  2660 => x"66c8799f",
  2661 => x"81eac149",
  2662 => x"c8799fc1",
  2663 => x"ecc14966",
  2664 => x"9fbf6e81",
  2665 => x"4966c879",
  2666 => x"c481eec1",
  2667 => x"799fbf66",
  2668 => x"c14966c8",
  2669 => x"9f6d81f0",
  2670 => x"cf4b7479",
  2671 => x"739bffff",
  2672 => x"4966c84a",
  2673 => x"7281f2c1",
  2674 => x"4a74799f",
  2675 => x"ffcf2ad0",
  2676 => x"4c729aff",
  2677 => x"c14966c8",
  2678 => x"9f7481f4",
  2679 => x"66c87379",
  2680 => x"81f8c149",
  2681 => x"72799f73",
  2682 => x"c14966c8",
  2683 => x"9f7281fa",
  2684 => x"268ee479",
  2685 => x"264c264d",
  2686 => x"694f264b",
  2687 => x"6953544d",
  2688 => x"696e694d",
  2689 => x"7267484d",
  2690 => x"6c646661",
  2691 => x"00652069",
  2692 => x"3030312e",
  2693 => x"20202020",
  2694 => x"69446500",
  2695 => x"6653544d",
  2696 => x"20792069",
  2697 => x"20202020",
  2698 => x"20202020",
  2699 => x"20202020",
  2700 => x"20202020",
  2701 => x"20202020",
  2702 => x"20202020",
  2703 => x"20202020",
  2704 => x"731e0020",
  2705 => x"d44b711e",
  2706 => x"87d40266",
  2707 => x"d84966c8",
  2708 => x"c84a7331",
  2709 => x"49a17232",
  2710 => x"718166cc",
  2711 => x"87e3c048",
  2712 => x"c24966d0",
  2713 => x"c6c491e8",
  2714 => x"dcc281d2",
  2715 => x"4a6a4aa1",
  2716 => x"66c89273",
  2717 => x"81e0c282",
  2718 => x"91724969",
  2719 => x"c18166cc",
  2720 => x"fd487189",
  2721 => x"711e87f1",
  2722 => x"49d4ff4a",
  2723 => x"c848d0ff",
  2724 => x"d0c278c5",
  2725 => x"7979c079",
  2726 => x"79797979",
  2727 => x"79727979",
  2728 => x"66c479c0",
  2729 => x"c879c079",
  2730 => x"79c07966",
  2731 => x"c07966cc",
  2732 => x"7966d079",
  2733 => x"66d479c0",
  2734 => x"2678c479",
  2735 => x"4a711e4f",
  2736 => x"9749a2c6",
  2737 => x"f0c34969",
  2738 => x"c01e7199",
  2739 => x"1ec11e1e",
  2740 => x"fe491ec0",
  2741 => x"d0c287f0",
  2742 => x"87f4f649",
  2743 => x"4f268eec",
  2744 => x"1e1ec01e",
  2745 => x"c11e1e1e",
  2746 => x"87dafe49",
  2747 => x"f649d0c2",
  2748 => x"8eec87de",
  2749 => x"711e4f26",
  2750 => x"48d0ff4a",
  2751 => x"ff78c5c8",
  2752 => x"e0c248d4",
  2753 => x"7878c078",
  2754 => x"c8787878",
  2755 => x"49721ec0",
  2756 => x"87e1d9fd",
  2757 => x"c448d0ff",
  2758 => x"4f262678",
  2759 => x"5c5b5e0e",
  2760 => x"86f80e5d",
  2761 => x"a2c24a71",
  2762 => x"7b97c14b",
  2763 => x"c14ca2c3",
  2764 => x"49a27c97",
  2765 => x"a2c451c0",
  2766 => x"7d97c04d",
  2767 => x"6e7ea2c5",
  2768 => x"c450c048",
  2769 => x"a2c648a6",
  2770 => x"4866c478",
  2771 => x"66d850c0",
  2772 => x"d2f0c31e",
  2773 => x"87eaf549",
  2774 => x"bf9766c8",
  2775 => x"66c81e49",
  2776 => x"1e49bf97",
  2777 => x"141e4915",
  2778 => x"49131e49",
  2779 => x"fc49c01e",
  2780 => x"49c887d4",
  2781 => x"c387d9f4",
  2782 => x"fd49d2f0",
  2783 => x"49d087f8",
  2784 => x"e087cdf4",
  2785 => x"87ebf98e",
  2786 => x"c64a711e",
  2787 => x"699749a2",
  2788 => x"a2c51e49",
  2789 => x"49699749",
  2790 => x"49a2c41e",
  2791 => x"1e496997",
  2792 => x"9749a2c3",
  2793 => x"c21e4969",
  2794 => x"699749a2",
  2795 => x"49c01e49",
  2796 => x"c287d3fb",
  2797 => x"d7f349d0",
  2798 => x"268eec87",
  2799 => x"1e731e4f",
  2800 => x"a2c24a71",
  2801 => x"d04b1149",
  2802 => x"c806abb7",
  2803 => x"49d1c287",
  2804 => x"d587fdf2",
  2805 => x"4966c887",
  2806 => x"c491e8c2",
  2807 => x"c281d2c6",
  2808 => x"797381e4",
  2809 => x"f249d0c2",
  2810 => x"caf887e6",
  2811 => x"1e731e87",
  2812 => x"a3c64b71",
  2813 => x"49699749",
  2814 => x"49a3c51e",
  2815 => x"1e496997",
  2816 => x"9749a3c4",
  2817 => x"c31e4969",
  2818 => x"699749a3",
  2819 => x"a3c21e49",
  2820 => x"49699749",
  2821 => x"4aa3c11e",
  2822 => x"e9f94912",
  2823 => x"49d0c287",
  2824 => x"ec87edf1",
  2825 => x"87cff78e",
  2826 => x"5c5b5e0e",
  2827 => x"711e0e5d",
  2828 => x"c2496e7e",
  2829 => x"7997c181",
  2830 => x"83c34b6e",
  2831 => x"6e7b97c1",
  2832 => x"c082c14a",
  2833 => x"4c6e7a97",
  2834 => x"97c084c4",
  2835 => x"c54d6e7c",
  2836 => x"6e55c085",
  2837 => x"9785c64d",
  2838 => x"c01e4d6d",
  2839 => x"4c6c971e",
  2840 => x"4b6b971e",
  2841 => x"4969971e",
  2842 => x"f849121e",
  2843 => x"d0c287d8",
  2844 => x"87dcf049",
  2845 => x"faf58ee8",
  2846 => x"5b5e0e87",
  2847 => x"ff0e5d5c",
  2848 => x"4c7186dc",
  2849 => x"1149a4c3",
  2850 => x"4aa4c44d",
  2851 => x"9749a4c5",
  2852 => x"31c84969",
  2853 => x"484a6a97",
  2854 => x"a6d4b071",
  2855 => x"7ea4c658",
  2856 => x"49bf976e",
  2857 => x"d898cf48",
  2858 => x"487158a6",
  2859 => x"dc98c0c1",
  2860 => x"ec4858a6",
  2861 => x"78a4c280",
  2862 => x"bf9766c4",
  2863 => x"c3059b4b",
  2864 => x"4bc0c487",
  2865 => x"c01e66d8",
  2866 => x"751e66f8",
  2867 => x"66e0c01e",
  2868 => x"66e0c01e",
  2869 => x"87eaf549",
  2870 => x"497086d0",
  2871 => x"59a6e0c0",
  2872 => x"c5029b73",
  2873 => x"f8c087fb",
  2874 => x"87c50266",
  2875 => x"c55ba6d0",
  2876 => x"48a6cc87",
  2877 => x"66cc78c1",
  2878 => x"66f8c04c",
  2879 => x"c087de02",
  2880 => x"c24966f4",
  2881 => x"c6c491e8",
  2882 => x"e4c281d2",
  2883 => x"48a6c881",
  2884 => x"66cc7869",
  2885 => x"b766c848",
  2886 => x"87c106a8",
  2887 => x"66fcc04c",
  2888 => x"c887d905",
  2889 => x"87e8ed49",
  2890 => x"7087fded",
  2891 => x"0599c449",
  2892 => x"f3ed87ca",
  2893 => x"c4497087",
  2894 => x"87f60299",
  2895 => x"88c14874",
  2896 => x"7058a6d0",
  2897 => x"029c744a",
  2898 => x"c187d4c1",
  2899 => x"c2c102ab",
  2900 => x"66f4c087",
  2901 => x"91e8c249",
  2902 => x"48d2c6c4",
  2903 => x"a6cc8071",
  2904 => x"4966c858",
  2905 => x"6981e0c2",
  2906 => x"e4c005ad",
  2907 => x"d44dc187",
  2908 => x"80c14866",
  2909 => x"c858a6d8",
  2910 => x"dcc24966",
  2911 => x"05a86981",
  2912 => x"a6d487d1",
  2913 => x"d078c048",
  2914 => x"80c14866",
  2915 => x"c258a6d4",
  2916 => x"c185c187",
  2917 => x"c149728b",
  2918 => x"0599718a",
  2919 => x"d887ecfe",
  2920 => x"87d90266",
  2921 => x"66dc4974",
  2922 => x"c34a7181",
  2923 => x"4d729aff",
  2924 => x"b7c84a71",
  2925 => x"5aa6d42a",
  2926 => x"a629b7d8",
  2927 => x"bf976e59",
  2928 => x"99f0c349",
  2929 => x"71b166d4",
  2930 => x"4966d41e",
  2931 => x"7129b7c8",
  2932 => x"1e66d81e",
  2933 => x"66d41e75",
  2934 => x"1e49bf97",
  2935 => x"e5f249c0",
  2936 => x"c086d487",
  2937 => x"c10566fc",
  2938 => x"49d087f1",
  2939 => x"c087e1ea",
  2940 => x"c24966f4",
  2941 => x"c6c491e8",
  2942 => x"807148d2",
  2943 => x"c858a6cc",
  2944 => x"81c84966",
  2945 => x"cdc10269",
  2946 => x"4966dc87",
  2947 => x"1e7131c9",
  2948 => x"fd4966cc",
  2949 => x"c487e7f5",
  2950 => x"a6e0c086",
  2951 => x"7866cc48",
  2952 => x"c0029c74",
  2953 => x"1ec087f5",
  2954 => x"fd4966cc",
  2955 => x"c187ddef",
  2956 => x"4966d01e",
  2957 => x"87f3edfd",
  2958 => x"66dc86c8",
  2959 => x"c080c148",
  2960 => x"c058a6e0",
  2961 => x"484966e0",
  2962 => x"e4c088c1",
  2963 => x"997158a6",
  2964 => x"87d2ff05",
  2965 => x"49c987c5",
  2966 => x"7387f5e8",
  2967 => x"c5fa059b",
  2968 => x"66fcc087",
  2969 => x"d087c502",
  2970 => x"87e4e849",
  2971 => x"ee8edcff",
  2972 => x"5e0e87c1",
  2973 => x"0e5d5c5b",
  2974 => x"4c7186e0",
  2975 => x"1149a4c3",
  2976 => x"58a6d448",
  2977 => x"c54aa4c4",
  2978 => x"699749a4",
  2979 => x"9731c849",
  2980 => x"71484a6a",
  2981 => x"58a6d8b0",
  2982 => x"6e7ea4c6",
  2983 => x"4d49bf97",
  2984 => x"48719dcf",
  2985 => x"dc98c0c1",
  2986 => x"ec4858a6",
  2987 => x"78a4c280",
  2988 => x"bf9766c4",
  2989 => x"1e66d84b",
  2990 => x"1e66f4c0",
  2991 => x"751e66d8",
  2992 => x"66e4c01e",
  2993 => x"87faed49",
  2994 => x"497086d0",
  2995 => x"59a6e0c0",
  2996 => x"c3059b73",
  2997 => x"4bc0c487",
  2998 => x"f3e649c4",
  2999 => x"4966dc87",
  3000 => x"1e7131c9",
  3001 => x"4966f4c0",
  3002 => x"c491e8c2",
  3003 => x"7148d2c6",
  3004 => x"58a6d480",
  3005 => x"fd4966d0",
  3006 => x"c487c3f2",
  3007 => x"029b7386",
  3008 => x"c087dfc4",
  3009 => x"c40266f4",
  3010 => x"c24a7387",
  3011 => x"724ac187",
  3012 => x"66f4c04c",
  3013 => x"cc87d302",
  3014 => x"e4c24966",
  3015 => x"48a6c881",
  3016 => x"66c87869",
  3017 => x"c106aab7",
  3018 => x"9c744c87",
  3019 => x"87d5c202",
  3020 => x"7087f5e5",
  3021 => x"0599c849",
  3022 => x"ebe587ca",
  3023 => x"c8497087",
  3024 => x"87f60299",
  3025 => x"c848d0ff",
  3026 => x"d4ff78c5",
  3027 => x"78f0c248",
  3028 => x"787878c0",
  3029 => x"c0c87878",
  3030 => x"d2f0c31e",
  3031 => x"eac8fd49",
  3032 => x"48d0ff87",
  3033 => x"f0c378c4",
  3034 => x"66d41ed2",
  3035 => x"deebfd49",
  3036 => x"d81ec187",
  3037 => x"e8fd4966",
  3038 => x"86cc87f1",
  3039 => x"c14866dc",
  3040 => x"a6e0c080",
  3041 => x"02abc158",
  3042 => x"cc87f3c0",
  3043 => x"e0c24966",
  3044 => x"4866d081",
  3045 => x"dd05a869",
  3046 => x"48a6d087",
  3047 => x"cc8578c1",
  3048 => x"dcc24966",
  3049 => x"05ad6981",
  3050 => x"4dc087d4",
  3051 => x"c14866d4",
  3052 => x"58a6d880",
  3053 => x"66d087c8",
  3054 => x"d480c148",
  3055 => x"8bc158a6",
  3056 => x"ebfd058c",
  3057 => x"0266d887",
  3058 => x"66dc87da",
  3059 => x"99ffc349",
  3060 => x"dc59a6d4",
  3061 => x"b7c84966",
  3062 => x"59a6d829",
  3063 => x"d84966dc",
  3064 => x"4d7129b7",
  3065 => x"49bf976e",
  3066 => x"7599f0c3",
  3067 => x"d81e71b1",
  3068 => x"b7c84966",
  3069 => x"dc1e7129",
  3070 => x"66dc1e66",
  3071 => x"9766d41e",
  3072 => x"c01e49bf",
  3073 => x"87fee949",
  3074 => x"9b7386d4",
  3075 => x"d087c702",
  3076 => x"87fce149",
  3077 => x"d0c287c6",
  3078 => x"87f4e149",
  3079 => x"fb059b73",
  3080 => x"8ee087e1",
  3081 => x"0e87cce7",
  3082 => x"5d5c5b5e",
  3083 => x"7186f80e",
  3084 => x"49a4c84c",
  3085 => x"2ac94a69",
  3086 => x"c3029a72",
  3087 => x"1e7287ca",
  3088 => x"4ad14972",
  3089 => x"87c8c3fd",
  3090 => x"99714a26",
  3091 => x"87c4c205",
  3092 => x"c0c0c4c1",
  3093 => x"fbc101aa",
  3094 => x"cc7ed187",
  3095 => x"01aac0f0",
  3096 => x"4dc487c5",
  3097 => x"7287ccc1",
  3098 => x"c649721e",
  3099 => x"dfc2fd4a",
  3100 => x"714a2687",
  3101 => x"87cc0599",
  3102 => x"aac0e0d9",
  3103 => x"c687c501",
  3104 => x"87efc04d",
  3105 => x"1e724bc5",
  3106 => x"4a734972",
  3107 => x"87c0c2fd",
  3108 => x"99714a26",
  3109 => x"7387cb05",
  3110 => x"c0d0c449",
  3111 => x"06aa7191",
  3112 => x"abc587cf",
  3113 => x"c187c205",
  3114 => x"d083c183",
  3115 => x"d5ff04ab",
  3116 => x"724d7387",
  3117 => x"7549721e",
  3118 => x"d3c1fd4a",
  3119 => x"26497087",
  3120 => x"721e714a",
  3121 => x"fd4ad11e",
  3122 => x"2687c5c1",
  3123 => x"c849264a",
  3124 => x"87db58a6",
  3125 => x"d07effc0",
  3126 => x"c449724d",
  3127 => x"721e7129",
  3128 => x"4affc01e",
  3129 => x"87e8c0fd",
  3130 => x"49264a26",
  3131 => x"c258a6c8",
  3132 => x"c449a4d8",
  3133 => x"dcc27966",
  3134 => x"797549a4",
  3135 => x"49a4e0c2",
  3136 => x"e4c2796e",
  3137 => x"79c149a4",
  3138 => x"e6e38ef8",
  3139 => x"49c01e87",
  3140 => x"bfdac6c4",
  3141 => x"c187c202",
  3142 => x"c2c9c449",
  3143 => x"87c202bf",
  3144 => x"d0ffb1c2",
  3145 => x"78c5c848",
  3146 => x"c348d4ff",
  3147 => x"787178fa",
  3148 => x"c448d0ff",
  3149 => x"1e4f2678",
  3150 => x"4a711e73",
  3151 => x"4966cc1e",
  3152 => x"c491e8c2",
  3153 => x"714bd2c6",
  3154 => x"fd497383",
  3155 => x"c487f0de",
  3156 => x"02987086",
  3157 => x"497387cb",
  3158 => x"87f5e7fd",
  3159 => x"c6fb4973",
  3160 => x"87e9fe87",
  3161 => x"0e87d0e2",
  3162 => x"5d5c5b5e",
  3163 => x"ff86f40e",
  3164 => x"7087f5dc",
  3165 => x"0299c449",
  3166 => x"ff87ecc5",
  3167 => x"c5c848d0",
  3168 => x"48d4ff78",
  3169 => x"c078c0c2",
  3170 => x"78787878",
  3171 => x"d4ff4d78",
  3172 => x"7678c048",
  3173 => x"ff49a54a",
  3174 => x"7997bfd4",
  3175 => x"c048d4ff",
  3176 => x"c1516878",
  3177 => x"adb7c885",
  3178 => x"ff87e304",
  3179 => x"78c448d0",
  3180 => x"486697c6",
  3181 => x"7058a6cc",
  3182 => x"c49bd04b",
  3183 => x"49732bb7",
  3184 => x"c491e8c2",
  3185 => x"c881d2c6",
  3186 => x"ca056981",
  3187 => x"49d1c287",
  3188 => x"87fcdaff",
  3189 => x"c787d0c4",
  3190 => x"494c6697",
  3191 => x"d099f0c3",
  3192 => x"87cc05a9",
  3193 => x"49721e73",
  3194 => x"c487d2e3",
  3195 => x"87f7c386",
  3196 => x"05acd0c2",
  3197 => x"497287c8",
  3198 => x"c387e5e3",
  3199 => x"ecc387e9",
  3200 => x"87ce05ac",
  3201 => x"1e731ec0",
  3202 => x"cfe44972",
  3203 => x"c386c887",
  3204 => x"d1c287d5",
  3205 => x"87cc05ac",
  3206 => x"49721e73",
  3207 => x"c487e9e5",
  3208 => x"87c3c386",
  3209 => x"05acc6c3",
  3210 => x"1e7387cc",
  3211 => x"cce64972",
  3212 => x"c286c487",
  3213 => x"e0c087f1",
  3214 => x"87cf05ac",
  3215 => x"731e1ec0",
  3216 => x"e849721e",
  3217 => x"86cc87f3",
  3218 => x"c387dcc2",
  3219 => x"d005acc4",
  3220 => x"c11ec087",
  3221 => x"721e731e",
  3222 => x"87dde849",
  3223 => x"c6c286cc",
  3224 => x"acf0c087",
  3225 => x"c087ce05",
  3226 => x"721e731e",
  3227 => x"87c2f049",
  3228 => x"f2c186c8",
  3229 => x"acc5c387",
  3230 => x"c187ce05",
  3231 => x"721e731e",
  3232 => x"87eeef49",
  3233 => x"dec186c8",
  3234 => x"05acc887",
  3235 => x"1e7387cc",
  3236 => x"d3e64972",
  3237 => x"c186c487",
  3238 => x"c0c187cd",
  3239 => x"87d005ac",
  3240 => x"1ec01ec1",
  3241 => x"49721e73",
  3242 => x"cc87cee7",
  3243 => x"87f7c086",
  3244 => x"cc059c74",
  3245 => x"721e7387",
  3246 => x"87f1e449",
  3247 => x"e6c086c4",
  3248 => x"1e66c887",
  3249 => x"496697c9",
  3250 => x"6697cc1e",
  3251 => x"97cf1e49",
  3252 => x"d21e4966",
  3253 => x"1e496697",
  3254 => x"deff49c4",
  3255 => x"86d487e8",
  3256 => x"ff49d1c2",
  3257 => x"f487e9d6",
  3258 => x"c6dcff8e",
  3259 => x"5b5e0e87",
  3260 => x"1e0e5d5c",
  3261 => x"d4ff7e71",
  3262 => x"c41e6e4b",
  3263 => x"fd49e2cb",
  3264 => x"c487fcd7",
  3265 => x"9d4d7086",
  3266 => x"87c3c302",
  3267 => x"bfeacbc4",
  3268 => x"fd496e4c",
  3269 => x"ff87cff4",
  3270 => x"c5c848d0",
  3271 => x"7bd6c178",
  3272 => x"7b154ac0",
  3273 => x"e0c082c1",
  3274 => x"f504aab7",
  3275 => x"48d0ff87",
  3276 => x"c5c878c4",
  3277 => x"7bd3c178",
  3278 => x"78c47bc1",
  3279 => x"c1029c74",
  3280 => x"f0c387fc",
  3281 => x"c0c87ed2",
  3282 => x"b7c08c4d",
  3283 => x"87c603ac",
  3284 => x"4da4c0c8",
  3285 => x"fdc34cc0",
  3286 => x"49bf97c3",
  3287 => x"d20299d0",
  3288 => x"c41ec087",
  3289 => x"fd49e2cb",
  3290 => x"c487e1da",
  3291 => x"4a497086",
  3292 => x"c387efc0",
  3293 => x"c41ed2f0",
  3294 => x"fd49e2cb",
  3295 => x"c487cdda",
  3296 => x"4a497086",
  3297 => x"c848d0ff",
  3298 => x"d4c178c5",
  3299 => x"bf976e7b",
  3300 => x"c1486e7b",
  3301 => x"c17e7080",
  3302 => x"f0ff058d",
  3303 => x"48d0ff87",
  3304 => x"9a7278c4",
  3305 => x"c087c505",
  3306 => x"87e5c048",
  3307 => x"cbc41ec1",
  3308 => x"d7fd49e2",
  3309 => x"86c487f5",
  3310 => x"fe059c74",
  3311 => x"d0ff87c4",
  3312 => x"78c5c848",
  3313 => x"c07bd3c1",
  3314 => x"c178c47b",
  3315 => x"c087c248",
  3316 => x"4d262648",
  3317 => x"4b264c26",
  3318 => x"1e004f26",
  3319 => x"bfc4d0c3",
  3320 => x"c3b9c149",
  3321 => x"ff59c8d0",
  3322 => x"ffc348d4",
  3323 => x"48d0ff78",
  3324 => x"ff78e1c8",
  3325 => x"78c148d4",
  3326 => x"787131c4",
  3327 => x"c048d0ff",
  3328 => x"4f2678e0",
  3329 => x"00000000",
  3330 => x"5c5b5e0e",
  3331 => x"4c711e0e",
  3332 => x"87ccfdfe",
  3333 => x"66d04b70",
  3334 => x"efc0c41e",
  3335 => x"e2dcfe49",
  3336 => x"7386c487",
  3337 => x"87d9059b",
  3338 => x"4aa4f4c0",
  3339 => x"49a4f0c0",
  3340 => x"66d08269",
  3341 => x"c1486952",
  3342 => x"6e7e7080",
  3343 => x"7098cf48",
  3344 => x"87c22679",
  3345 => x"4c264d26",
  3346 => x"4f264b26",
  3347 => x"5c5b5e0e",
  3348 => x"cc4b710e",
  3349 => x"c2494c66",
  3350 => x"ca0299c0",
  3351 => x"1ee0c387",
  3352 => x"e3fe4973",
  3353 => x"7486c487",
  3354 => x"99c0c449",
  3355 => x"c287c502",
  3356 => x"87c3b4c0",
  3357 => x"749cffc1",
  3358 => x"fe49731e",
  3359 => x"ff2687ca",
  3360 => x"731e87c4",
  3361 => x"d3c31e1e",
  3362 => x"ff49bfe8",
  3363 => x"7087c8c8",
  3364 => x"cfc10298",
  3365 => x"e6cec487",
  3366 => x"cec448bf",
  3367 => x"02a8bfea",
  3368 => x"c487c1c1",
  3369 => x"c44beece",
  3370 => x"83bfe6ce",
  3371 => x"c04b6b97",
  3372 => x"c7ff49e8",
  3373 => x"497087d5",
  3374 => x"59ecd3c3",
  3375 => x"c848d0ff",
  3376 => x"d4ff78e1",
  3377 => x"7378c548",
  3378 => x"08d4ff48",
  3379 => x"48d0ff78",
  3380 => x"c478e0c0",
  3381 => x"48bfe6ce",
  3382 => x"7e7080c1",
  3383 => x"98cf486e",
  3384 => x"58eacec4",
  3385 => x"87e0fd26",
  3386 => x"00000000",
  3387 => x"5c5b5e0e",
  3388 => x"d8ff0e5d",
  3389 => x"c47ec086",
  3390 => x"49bffecd",
  3391 => x"1e7181c2",
  3392 => x"4ac61e72",
  3393 => x"87fcf0fc",
  3394 => x"4a264871",
  3395 => x"a6c84926",
  3396 => x"fecdc458",
  3397 => x"81c449bf",
  3398 => x"1e721e71",
  3399 => x"f0fc4ac6",
  3400 => x"487187e2",
  3401 => x"49264a26",
  3402 => x"fd58a6cc",
  3403 => x"dfc387d4",
  3404 => x"ff49bff6",
  3405 => x"7087e0c5",
  3406 => x"f3ca0298",
  3407 => x"ff49d087",
  3408 => x"7087c8c5",
  3409 => x"fadfc349",
  3410 => x"744cc059",
  3411 => x"fe91c449",
  3412 => x"4a6981d0",
  3413 => x"cdc44974",
  3414 => x"c481bffe",
  3415 => x"cecec491",
  3416 => x"9a797281",
  3417 => x"7287d202",
  3418 => x"7189c149",
  3419 => x"c1486e9a",
  3420 => x"727e7080",
  3421 => x"eeff059a",
  3422 => x"c284c187",
  3423 => x"ff04acb7",
  3424 => x"486e87c9",
  3425 => x"a8b7fcc0",
  3426 => x"87e4c904",
  3427 => x"4a744cc0",
  3428 => x"c48266c4",
  3429 => x"cecec492",
  3430 => x"c8497482",
  3431 => x"91c48166",
  3432 => x"81cecec4",
  3433 => x"49694a6a",
  3434 => x"4b74b972",
  3435 => x"bffecdc4",
  3436 => x"c493c483",
  3437 => x"6b83cece",
  3438 => x"714872ba",
  3439 => x"58a6d498",
  3440 => x"cdc44974",
  3441 => x"c481bffe",
  3442 => x"cecec491",
  3443 => x"d47e6981",
  3444 => x"78c048a6",
  3445 => x"c35ca6d0",
  3446 => x"66d04cff",
  3447 => x"0229df49",
  3448 => x"cc87dcc7",
  3449 => x"e0c04a66",
  3450 => x"8266d492",
  3451 => x"7248ffc0",
  3452 => x"d84a7088",
  3453 => x"78c048a6",
  3454 => x"78c080c4",
  3455 => x"29df496e",
  3456 => x"59a6e4c0",
  3457 => x"48facdc4",
  3458 => x"497278c1",
  3459 => x"2ab731c3",
  3460 => x"ffc0b172",
  3461 => x"c391c499",
  3462 => x"714deceb",
  3463 => x"494b6d85",
  3464 => x"99c0c0c4",
  3465 => x"c087d702",
  3466 => x"c00266e0",
  3467 => x"80c887c7",
  3468 => x"cac678c0",
  3469 => x"c2cec487",
  3470 => x"c678c148",
  3471 => x"e0c087c1",
  3472 => x"87d80266",
  3473 => x"c0c24973",
  3474 => x"c00299c0",
  3475 => x"b7d087c3",
  3476 => x"fd486d2b",
  3477 => x"7098ffff",
  3478 => x"87fac07d",
  3479 => x"bfc2cec4",
  3480 => x"87f2c002",
  3481 => x"b7d04873",
  3482 => x"a6e8c028",
  3483 => x"02987058",
  3484 => x"c487e3c0",
  3485 => x"49bfcace",
  3486 => x"99c0e0c0",
  3487 => x"87cac002",
  3488 => x"e0c04970",
  3489 => x"c00299c0",
  3490 => x"486d87cc",
  3491 => x"b0c0c0c2",
  3492 => x"e4c07d70",
  3493 => x"49734b66",
  3494 => x"99c0c0c8",
  3495 => x"87ffc202",
  3496 => x"0266e0c0",
  3497 => x"7387c8c0",
  3498 => x"9ac0cc4a",
  3499 => x"f387cfc0",
  3500 => x"cec49bff",
  3501 => x"cc4abfca",
  3502 => x"b3729ac0",
  3503 => x"9a727d73",
  3504 => x"4887df02",
  3505 => x"c088c0c4",
  3506 => x"7058a6e8",
  3507 => x"e0c00298",
  3508 => x"c0c44887",
  3509 => x"a6e8c088",
  3510 => x"02987058",
  3511 => x"c187c2c1",
  3512 => x"497387ef",
  3513 => x"91c29974",
  3514 => x"81e0ebc3",
  3515 => x"eec14b11",
  3516 => x"74497387",
  3517 => x"c391c299",
  3518 => x"c181e0eb",
  3519 => x"c44b1181",
  3520 => x"49bfcace",
  3521 => x"c099c0c4",
  3522 => x"029966e0",
  3523 => x"dc87c9c0",
  3524 => x"eac048a6",
  3525 => x"87c7c178",
  3526 => x"c448a6d8",
  3527 => x"fec078ea",
  3528 => x"74497387",
  3529 => x"c391c299",
  3530 => x"c181e0eb",
  3531 => x"c44b1181",
  3532 => x"49bfcace",
  3533 => x"c099c0c8",
  3534 => x"029966e0",
  3535 => x"dc87c9c0",
  3536 => x"f6c048a6",
  3537 => x"87d7c078",
  3538 => x"c448a6d8",
  3539 => x"cec078f6",
  3540 => x"74497387",
  3541 => x"c391c299",
  3542 => x"c181e0eb",
  3543 => x"c04b1181",
  3544 => x"c00266e0",
  3545 => x"497387db",
  3546 => x"fcc7b9ff",
  3547 => x"487199c0",
  3548 => x"bfcacec4",
  3549 => x"cecec498",
  3550 => x"c49b7458",
  3551 => x"d3c0b3c0",
  3552 => x"c7497387",
  3553 => x"7199c0fc",
  3554 => x"cacec448",
  3555 => x"cec4b0bf",
  3556 => x"9b7458ce",
  3557 => x"c00266d8",
  3558 => x"c41e87ca",
  3559 => x"f249facd",
  3560 => x"86c487ea",
  3561 => x"cdc41e73",
  3562 => x"dff249fa",
  3563 => x"dc86c487",
  3564 => x"cac00266",
  3565 => x"cdc41e87",
  3566 => x"cff249fa",
  3567 => x"d086c487",
  3568 => x"30c14866",
  3569 => x"6e58a6d4",
  3570 => x"7030c148",
  3571 => x"4866d47e",
  3572 => x"a6d880c1",
  3573 => x"b7e0c058",
  3574 => x"fdf704a8",
  3575 => x"4c66cc87",
  3576 => x"b7c284c1",
  3577 => x"e5f604ac",
  3578 => x"fecdc487",
  3579 => x"7866c448",
  3580 => x"f18ed8ff",
  3581 => x"000087ce",
  3582 => x"c01e0000",
  3583 => x"c449724a",
  3584 => x"cecec491",
  3585 => x"c179ff81",
  3586 => x"aab7c682",
  3587 => x"c487ee04",
  3588 => x"c048fecd",
  3589 => x"80c87840",
  3590 => x"4f2678c0",
  3591 => x"711e731e",
  3592 => x"87c8f34b",
  3593 => x"d0fe4973",
  3594 => x"dbf087ca",
  3595 => x"5b5e0e87",
  3596 => x"711e0e5c",
  3597 => x"d04bc04c",
  3598 => x"e9c00266",
  3599 => x"8ac14a87",
  3600 => x"87e2c002",
  3601 => x"87de028a",
  3602 => x"028aeec0",
  3603 => x"c187c6c1",
  3604 => x"727e738a",
  3605 => x"d7c1029a",
  3606 => x"738ac187",
  3607 => x"029a727e",
  3608 => x"c187cdc1",
  3609 => x"9c7487d9",
  3610 => x"87d3c102",
  3611 => x"c1026c97",
  3612 => x"c0c487cd",
  3613 => x"c148bff9",
  3614 => x"fdc0c4b0",
  3615 => x"c0d6fe58",
  3616 => x"4966d087",
  3617 => x"cfc381c1",
  3618 => x"745997de",
  3619 => x"87dde949",
  3620 => x"eac04b70",
  3621 => x"4b66d087",
  3622 => x"738bf0c0",
  3623 => x"fe49c01e",
  3624 => x"7387ebfd",
  3625 => x"fe49741e",
  3626 => x"c887e3fd",
  3627 => x"87e0c086",
  3628 => x"c04966d0",
  3629 => x"1e7189f1",
  3630 => x"fae14974",
  3631 => x"c486c487",
  3632 => x"48bff9c0",
  3633 => x"c0c498fe",
  3634 => x"d4fe58fd",
  3635 => x"487387f3",
  3636 => x"87f2ed26",
  3637 => x"c01e731e",
  3638 => x"f9c0c44b",
  3639 => x"b0c148bf",
  3640 => x"58fdc0c4",
  3641 => x"87d9d4fe",
  3642 => x"48ccc4c1",
  3643 => x"1ec850c0",
  3644 => x"49fecec4",
  3645 => x"87eddbfd",
  3646 => x"1e7286c4",
  3647 => x"48dce6c3",
  3648 => x"49c6cfc4",
  3649 => x"204aa1c4",
  3650 => x"05aa7141",
  3651 => x"4a2687f9",
  3652 => x"49fecec4",
  3653 => x"87c6fefc",
  3654 => x"029a4a70",
  3655 => x"fd4987c5",
  3656 => x"7287f5ce",
  3657 => x"e0e6c31e",
  3658 => x"c6cfc448",
  3659 => x"4aa1c449",
  3660 => x"aa714120",
  3661 => x"87f8ff05",
  3662 => x"1ec04a26",
  3663 => x"49fecec4",
  3664 => x"87cafbfe",
  3665 => x"1e7286c4",
  3666 => x"48e4e6c3",
  3667 => x"49c6cfc4",
  3668 => x"204aa1c4",
  3669 => x"05aa7141",
  3670 => x"2687f8ff",
  3671 => x"fecec44a",
  3672 => x"87c9e649",
  3673 => x"c0059870",
  3674 => x"e6c387c4",
  3675 => x"49c04be8",
  3676 => x"87c6ccfd",
  3677 => x"7387c3fa",
  3678 => x"c5c0029b",
  3679 => x"dbfc4987",
  3680 => x"49ca87e7",
  3681 => x"87c7dbfc",
  3682 => x"bff9c0c4",
  3683 => x"c498fe48",
  3684 => x"fe58fdc0",
  3685 => x"7387ead1",
  3686 => x"87ecea48",
  3687 => x"00202020",
  3688 => x"00444856",
  3689 => x"004d4f52",
  3690 => x"204d4f52",
  3691 => x"64616f6c",
  3692 => x"20676e69",
  3693 => x"6c696166",
  3694 => x"0e006465",
  3695 => x"5d5c5b5e",
  3696 => x"d7c11e0e",
  3697 => x"87f2f84d",
  3698 => x"fe87e1ec",
  3699 => x"fe87e9e9",
  3700 => x"ff87d1f5",
  3701 => x"6e87d0de",
  3702 => x"ffffc149",
  3703 => x"c1486e99",
  3704 => x"717e7080",
  3705 => x"87ca0599",
  3706 => x"87e9fdfd",
  3707 => x"cffe4970",
  3708 => x"497587e3",
  3709 => x"87c2ccfe",
  3710 => x"c24b4970",
  3711 => x"fe49dd9b",
  3712 => x"7087f7cb",
  3713 => x"fffe0298",
  3714 => x"029b7387",
  3715 => x"7587f9fe",
  3716 => x"e5cbfe49",
  3717 => x"05987087",
  3718 => x"49dd87cb",
  3719 => x"87dacbfe",
  3720 => x"de029870",
  3721 => x"fe49c187",
  3722 => x"7587c9c8",
  3723 => x"c9cbfe49",
  3724 => x"05987087",
  3725 => x"dd87eeff",
  3726 => x"fdcafe49",
  3727 => x"05987087",
  3728 => x"cf87e2ff",
  3729 => x"f1fe49e8",
  3730 => x"4b7087c1",
  3731 => x"ebc31ec0",
  3732 => x"effe49c9",
  3733 => x"86c487d8",
  3734 => x"fe494c73",
  3735 => x"7087f8f0",
  3736 => x"87cc0598",
  3737 => x"f0fe4974",
  3738 => x"987087ed",
  3739 => x"87f4ff02",
  3740 => x"e2fe49c0",
  3741 => x"497587f0",
  3742 => x"87fec9fe",
  3743 => x"99c24970",
  3744 => x"c187d405",
  3745 => x"ebc6fe49",
  3746 => x"fe497587",
  3747 => x"7087ebc9",
  3748 => x"0299c249",
  3749 => x"7587ecff",
  3750 => x"ddc9fe49",
  3751 => x"02987087",
  3752 => x"c187d2c0",
  3753 => x"cbc6fe49",
  3754 => x"fe497587",
  3755 => x"7087cbc9",
  3756 => x"eeff0598",
  3757 => x"1ee8cf87",
  3758 => x"49d3ebc3",
  3759 => x"87eeedfe",
  3760 => x"c3fc86c4",
  3761 => x"fbe52687",
  3762 => x"75615087",
  3763 => x"676e6973",
  3764 => x"55002e2e",
  3765 => x"7561706e",
  3766 => x"676e6973",
  3767 => x"002e2e2e",
  3768 => x"c8d0cbcd",
  3769 => x"3e3d3c3b",
  3770 => x"4241403f",
  3771 => x"00d2000e",
  3772 => x"009c001c",
  3773 => x"089d8000",
  3774 => x"00588005",
  3775 => x"00438002",
  3776 => x"00448003",
  3777 => x"00578004",
  3778 => x"08b88001",
  3779 => x"00000004",
  3780 => x"00000011",
  3781 => x"0000001e",
  3782 => x"00000005",
  3783 => x"0000002c",
  3784 => x"0000001f",
  3785 => x"00000012",
  3786 => x"0000012a",
  3787 => x"00000006",
  3788 => x"00000013",
  3789 => x"00000020",
  3790 => x"00000007",
  3791 => x"0000002e",
  3792 => x"00000021",
  3793 => x"00000014",
  3794 => x"0000002d",
  3795 => x"00470008",
  3796 => x"00000015",
  3797 => x"00000022",
  3798 => x"00480009",
  3799 => x"00000030",
  3800 => x"00000023",
  3801 => x"004b0016",
  3802 => x"0000002f",
  3803 => x"0049000a",
  3804 => x"004c0017",
  3805 => x"004f0024",
  3806 => x"00b5000b",
  3807 => x"00520032",
  3808 => x"00500025",
  3809 => x"004d0018",
  3810 => x"00000031",
  3811 => x"0000000d",
  3812 => x"00370019",
  3813 => x"00510026",
  3814 => x"0000000c",
  3815 => x"00530034",
  3816 => x"004a0027",
  3817 => x"0045001a",
  3818 => x"00000033",
  3819 => x"00cf0042",
  3820 => x"0037001b",
  3821 => x"00000028",
  3822 => x"00c700d3",
  3823 => x"00000236",
  3824 => x"002b0029",
  3825 => x"0000002b",
  3826 => x"004e0035",
  3827 => x"00450002",
  3828 => x"00580001",
  3829 => x"000f041d",
  3830 => x"00000003",
  3831 => x"00000039",
  3832 => x"00000038",
  3833 => x"00000010",
  3834 => x"00004000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
